// Seed: 561102826984812543,5224943229413370507

module vu
  ( output logic [4:1][0:3][1:2][4:3]  a
  , output shortint bifyijlrnu [3:3]
  , input supply1 logic [0:2] byt [2:2][2:1]
  , input wor logic [0:4][1:3][1:3] wej [4:2]
  , input wire logic [3:2][4:3][3:2] pziwea [3:2][2:3][4:3][3:0]
  , input logic [0:0][4:4][4:4] trxbyhw [2:3]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign byt = byt;
  assign pziwea = pziwea;
endmodule: vu

module bjwsy
  (output logic oheto [1:3], output supply0 logic czmgpod [1:0][3:0][2:1][2:2], input bit [2:0][2:4][3:4] umtmuyxnu [2:4]);
  
  
  and ev(anhfw, anhfw, fttjsglz);
  
  
  // Single-driven assigns
  assign oheto = '{'bx1,'b011,'b00001};
  
  // Multi-driven assigns
  assign fttjsglz = 'bx;
endmodule: bjwsy

module eaa
  (input uwire logic vsbr [4:3][2:2]);
  
  logic cunw [1:3];
  supply0 logic bmvxpfjq [1:0][3:0][2:1][2:2];
  logic yiwcotvx [1:3];
  bit [2:0][2:4][3:4] mtrtc [2:4];
  
  bjwsy ly(.oheto(yiwcotvx), .czmgpod(bmvxpfjq), .umtmuyxnu(mtrtc));
  
  bjwsy hfvibuzmer(.oheto(cunw), .czmgpod(bmvxpfjq), .umtmuyxnu(mtrtc));
  
  
  // Single-driven assigns
  assign mtrtc = mtrtc;
  
  // Multi-driven assigns
  assign bmvxpfjq = '{'{'{'{'b1},'{'bx}},'{'{'b0z},'{'bxz111}},'{'{'bz1x},'{'bx001}},'{'{'b11z},'{'b10x}}},'{'{'{'b00x},'{'b1}},'{'{'b01zz0},'{'bzxz0}},'{'{'b1z},'{'bx}},'{'{'b1010},'{'bx}}}};
endmodule: eaa



// Seed after: 2901206930565052048,5224943229413370507
