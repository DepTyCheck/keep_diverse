// Seed: 12814626189442541259,5224943229413370507

module xnbgo
  ( output realtime rrb
  , output reg [0:2]  rddteeresy
  , output logic [1:1]  mpgtznafr
  , output wand logic [0:4][4:1][1:3]  vcvzx
  , input reg [4:4][2:0] zr [2:2]
  , input tri0 logic nqp
  , input bit [1:0] eozwjhk [3:1][1:4][3:3]
  , input byte hzpiycocz
  );
  
  
  not zwy(umgb, rrb);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime rrb -> logic rrb
  
  or gmhyfu(d, rddteeresy, rrb);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2]  rddteeresy -> logic rddteeresy
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime rrb -> logic rrb
  
  or oqhnzjag(rrb, nqp, hzpiycocz);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic rrb -> realtime rrb
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte hzpiycocz -> logic hzpiycocz
  
  
  // Single-driven assigns
  assign rddteeresy = hzpiycocz;
  assign mpgtznafr = d;
  
  // Multi-driven assigns
endmodule: xnbgo

module gxmlkxl
  (output tri1 logic [3:2][1:2][2:2] wjad [2:0][2:1][4:4][3:4], input shortreal piohpebqy);
  
  bit [1:0] xsrjalsj [3:1][1:4][3:3];
  reg [4:4][2:0] sgnpyf [2:2];
  
  xnbgo m( .rrb(astspfvps)
         , .rddteeresy(k)
         , .mpgtznafr(jmncuq)
         , .vcvzx(uljobwxp)
         , .zr(sgnpyf)
         , .nqp(piohpebqy)
         , .eozwjhk(xsrjalsj)
         , .hzpiycocz(uljobwxp)
         );
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime rrb -> wire logic astspfvps
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2]  rddteeresy -> wire logic k
  //
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   wand logic [0:4][4:1][1:3]  vcvzx -> wire logic uljobwxp
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal piohpebqy -> tri0 logic nqp
  //
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic uljobwxp -> byte hzpiycocz
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign wjad = wjad;
  assign k = piohpebqy;
  assign uljobwxp = 'b00x;
endmodule: gxmlkxl



// Seed after: 4214566392895304490,5224943229413370507
