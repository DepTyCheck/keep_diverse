// Seed: 12148350361508476340,5224943229413370507

module h
  ( output uwire logic [3:1][4:4][2:4] rabefg [4:1][2:4]
  , output trireg logic [2:4][3:3][2:2][0:3] jyrxngbp [0:4][4:4]
  , output logic pbh
  , output supply1 logic [1:0][1:0]  aj
  , input triand logic uszcgau [4:3][4:0][0:2]
  );
  
  
  not toqzxmr(pbh, yda);
  
  
  // Single-driven assigns
  assign rabefg = rabefg;
  
  // Multi-driven assigns
  assign aj = pbh;
  assign jyrxngbp = jyrxngbp;
  assign yda = 'bx0xx0;
endmodule: h

module fzvwkztuz
  ( output shortreal ssylzac
  , output tri1 logic [4:2][1:4][1:3] mdtar [4:2][4:1]
  , output shortreal qbnq
  , input reg [0:2]  sbvkqk
  , input tri0 logic xzstxn [4:2][0:1][0:1][0:2]
  );
  
  
  and kqx(ssylzac, qbnq, ssylzac);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic ssylzac -> shortreal ssylzac
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal qbnq -> logic qbnq
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal ssylzac -> logic ssylzac
  
  
  // Single-driven assigns
  assign qbnq = 'bz0;
  
  // Multi-driven assigns
endmodule: fzvwkztuz



// Seed after: 3814454678116103976,5224943229413370507
