// Seed: 14781989141431543639,5224943229413370507

module bnfuknwiy
  (output reg xqyckrgv, output uwire logic [0:0]  gbtgbdv);
  
  
  and maja(xqyckrgv, xqyckrgv, pfpbylo);
  
  xor gl(mrik, wmp, xqyckrgv);
  
  and kvqrwcvqg(ukrlj, mkw, ukrlj);
  
  
  // Single-driven assigns
  assign gbtgbdv = gbtgbdv;
  
  // Multi-driven assigns
  assign wmp = 'bzz;
endmodule: bnfuknwiy

module kxe
  ( output uwire logic [4:1][3:0] etwlaiba [1:1][3:2]
  , output supply1 logic a [2:1][4:0][4:0]
  , input logic futa [0:4]
  , input bit [4:3]  peo
  );
  
  
  not rpxjluy(yankslkev, yankslkev);
  
  not r(yankslkev, tlhnexcv);
  
  xor wjab(yankslkev, yankslkev, yankslkev);
  
  bnfuknwiy cqdrwh(.xqyckrgv(spgjne), .gbtgbdv(vcirfiurb));
  
  
  // Single-driven assigns
  assign etwlaiba = etwlaiba;
  
  // Multi-driven assigns
endmodule: kxe

module jsahtm
  (output bit [3:1] tigfpszquy [0:0][2:2], output tri logic [1:2] chddbq [4:3][4:3][3:1][0:4]);
  
  uwire logic [4:1][3:0] yaxlbu [1:1][3:2];
  supply1 logic m [2:1][4:0][4:0];
  uwire logic [4:1][3:0] dkcrkzvzzs [1:1][3:2];
  logic zhapcshe [0:4];
  
  and iqnzl(he, he, fmmw);
  
  kxe c(.etwlaiba(dkcrkzvzzs), .a(m), .futa(zhapcshe), .peo(he));
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic he -> bit [4:3]  peo
  
  kxe yialwutu(.etwlaiba(yaxlbu), .a(m), .futa(zhapcshe), .peo(he));
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic he -> bit [4:3]  peo
  
  
  // Single-driven assigns
  assign tigfpszquy = '{'{'{'b00,'b11100,'b01101}}};
  assign zhapcshe = '{'bxx,'bz01,'b001,'bxx0x1,'bx};
  
  // Multi-driven assigns
  assign fmmw = he;
endmodule: jsahtm

module sear
  (output real yrcefobnb [1:1], output reg [1:2][0:0]  gly, output bit [0:4][3:3] ht [1:1], output wand logic [0:3]  yqgzzup);
  
  supply1 logic juioutypoj [2:1][4:0][4:0];
  uwire logic [4:1][3:0] vpsefyyn [1:1][3:2];
  logic wud [0:4];
  
  not uslsu(vkpjrp, botdsaekn);
  
  kxe rwzqpctayp(.etwlaiba(vpsefyyn), .a(juioutypoj), .futa(wud), .peo(lofqwmqjem));
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic lofqwmqjem -> bit [4:3]  peo
  
  or pvrondrgkw(gly, mvlwkm, lcrmkuy);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic gly -> reg [1:2][0:0]  gly
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign lcrmkuy = mvlwkm;
  assign lofqwmqjem = gly;
  assign botdsaekn = vkpjrp;
  assign yqgzzup = '{'b001,'bz,'bz0,'bz1};
  assign juioutypoj = '{'{'{'bx,'bz0zx0,'bxx1z,'b1,'b1x11x},'{'bx,'bxxzx0,'bxz0,'b1,'b11x},'{'bxx,'bxzx,'bx00,'b00,'bx},'{'bzx101,'b10,'b1xz,'bx0,'b1},'{'bz10xz,'b10,'bzz,'b0z,'b0z}},'{'{'bzzx1,'b1011,'b10,'b01x0z,'bxzx},'{'b1,'b1xz0,'bzz,'bxx,'bx1},'{'bx1x,'bz00x,'b10x00,'b0z01x,'bx001},'{'b011x1,'b00z0,'bz11zx,'bz01,'bzxx},'{'b0z010,'bz11,'b1xzz,'b011,'b0xz}}};
endmodule: sear



// Seed after: 5139529512849536609,5224943229413370507
