// Seed: 4993766961193060316,5224943229413370507

module ghwjqlqif
  ();
  
  
  not cvdda(ha, mk);
  
  xor fjju(wlwue, qah, zdyi);
  
  not dhg(wlwue, ha);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign mk = 'b0;
endmodule: ghwjqlqif

module ohyucut
  ( output shortreal xabcbgeij
  , input tri1 logic [2:3][1:4][3:3] nek [2:1][4:2][2:2][0:0]
  , input trireg logic [0:0][3:4][1:3] wudx [0:4][4:4][0:4]
  );
  
  
  not iupksx(pps, zakrobb);
  
  xor egvdzbi(epo, sthzgjjrh, xabcbgeij);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal xabcbgeij -> logic xabcbgeij
  
  or iwenlkfmmx(zfya, ljsclb, dcmeklu);
  
  
  // Single-driven assigns
  assign xabcbgeij = xabcbgeij;
  
  // Multi-driven assigns
  assign zakrobb = dcmeklu;
endmodule: ohyucut

module nqksnslgdt
  ( output supply1 logic [0:0][0:0][4:0]  axiue
  , output shortint e [3:4][4:4]
  , input wire logic [4:3][3:0] sgnew [3:3][1:0][4:3][2:4]
  , input logic cihs [2:1][4:4]
  );
  
  
  and v(axiue, unepkijwa, oxuptc);
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   logic axiue -> supply1 logic [0:0][0:0][4:0]  axiue
  
  or xsea(j, axiue, oxuptc);
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   supply1 logic [0:0][0:0][4:0]  axiue -> logic axiue
  
  or punr(axiue, rlfhkevoeb, uirvypva);
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   logic axiue -> supply1 logic [0:0][0:0][4:0]  axiue
  
  ghwjqlqif vaxube();
  
  
  // Single-driven assigns
  assign e = e;
  
  // Multi-driven assigns
  assign j = oxuptc;
endmodule: nqksnslgdt

module mftutjpyta
  ( output bit [4:0][4:0] hziez [4:0]
  , output triand logic [0:4][1:0] uuyzobx [1:1]
  , output trior logic [3:2][0:2] lvmixv [2:0]
  , output reg ixjpzpb [2:2][2:1]
  , input logic [3:1][1:2][2:0][4:2]  evrivbbdlj
  , input supply1 logic umff [4:0][1:1]
  );
  
  
  or qtkurl(otwhp, otwhp, otwhp);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: mftutjpyta



// Seed after: 9772030656613686378,5224943229413370507
