// Seed: 14061539277969093024,5224943229413370507

module svc
  ( output byte ajfnhbffii
  , output time neqc
  , output tri logic [2:4][3:1][2:1][3:0] ddhntxfl [1:3][0:2][4:3][3:3]
  , input tri1 logic [1:4][1:4][4:3] h [2:4][1:4][4:0][2:2]
  , input logic iluh
  , input shortint ioeuax [0:0]
  );
  
  
  not jlkif(neqc, neqc);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  //   logic neqc -> time neqc
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  //   time neqc -> logic neqc
  
  or c(m, ajfnhbffii, ajfnhbffii);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte ajfnhbffii -> logic ajfnhbffii
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte ajfnhbffii -> logic ajfnhbffii
  
  
  // Single-driven assigns
  assign ajfnhbffii = 'b0101;
  
  // Multi-driven assigns
  assign h = h;
  assign m = 'bx0z0;
  assign ddhntxfl = ddhntxfl;
endmodule: svc

module um
  ( output reg [0:2][2:2]  gnmhzkgc
  , output time wglrv
  , output integer mpdxupjbp [4:2]
  , input trior logic [3:0][3:4][2:0][1:1] nyci [0:4]
  , input logic jmmgqrga
  );
  
  
  or yrwivnye(btci, dmaft, gnmhzkgc);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][2:2]  gnmhzkgc -> logic gnmhzkgc
  
  
  // Single-driven assigns
  assign gnmhzkgc = '{'{'bx10},'{'bx},'{'bx}};
  assign mpdxupjbp = mpdxupjbp;
  assign wglrv = wglrv;
  
  // Multi-driven assigns
endmodule: um

module bnendouhcq
  ( output wand logic [3:2][1:4][4:4] xajepuf [3:4][1:0][2:1][0:2]
  , input tri1 logic [2:0] haypqz [1:2][4:1]
  , input reg [2:0][3:0] ynjoyfqj [1:4][1:0]
  , input logic gqogq
  , input shortreal wksoziudt [3:0]
  );
  
  integer ioqz [4:2];
  trior logic [3:0][3:4][2:0][1:1] zd [0:4];
  
  xor pfixvw(scawezub, gqogq, ig);
  
  um vwaukzzk(.gnmhzkgc(zqyuypbutm), .wglrv(szqzxpxa), .mpdxupjbp(ioqz), .nyci(zd), .jmmgqrga(gqogq));
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][2:2]  gnmhzkgc -> wire logic zqyuypbutm
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  //   time wglrv -> wire logic szqzxpxa
  
  and elfpvafomq(ig, zqvm, ig);
  
  not ytwedumvmd(nkzkdgwlgt, ztsdog);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xajepuf = xajepuf;
  assign zqyuypbutm = 'bxx0x0;
  assign zd = zd;
  assign ig = 'bz;
  assign haypqz = '{'{'{'bx,'bz00x1,'b00zx1},'{'bz0xxz,'bx11z,'b1011z},'{'b01x,'bxzx11,'bz0},'{'b0z,'b010x,'b101x}},'{'{'b0,'b0,'b110},'{'b0zzx,'bx00,'b11z00},'{'b1,'b0x,'b10x11},'{'b0x,'b11zz,'b1}}};
endmodule: bnendouhcq

module sejkvceskl
  (output logic pojm, output supply1 logic [0:0][3:4][2:1][2:3] clynhqy [1:0][3:0][3:4]);
  
  integer zwuy [4:2];
  trior logic [3:0][3:4][2:0][1:1] ykp [0:4];
  
  um xcal(.gnmhzkgc(pojm), .wglrv(l), .mpdxupjbp(zwuy), .nyci(ykp), .jmmgqrga(pojm));
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [0:2][2:2]  gnmhzkgc -> logic pojm
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  //   time wglrv -> wire logic l
  
  not gxdkzgc(l, pojm);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ykp = ykp;
  assign l = 'bz11;
  assign clynhqy = clynhqy;
endmodule: sejkvceskl



// Seed after: 5054388276277724192,5224943229413370507
