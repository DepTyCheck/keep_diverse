// Seed: 11869620239679120121,5224943229413370507

module dlcuctbxm
  (output tri0 logic [0:0][1:0] betoddf [4:0][3:3], output logic lfsopwxfyx [3:2], output tri1 logic [1:1][1:1] sgelmab [0:1][1:1]);
  
  
  not qf(omi, cxmqpotm);
  
  
  // Single-driven assigns
  assign lfsopwxfyx = '{'b1,'b0z};
  
  // Multi-driven assigns
  assign omi = cxmqpotm;
  assign sgelmab = sgelmab;
  assign betoddf = '{'{'{'{'b0xxx,'bz0xzx}}},'{'{'{'b1011z,'b10x1}}},'{'{'{'b101,'b0}}},'{'{'{'b0010,'b1zz}}},'{'{'{'b0,'b00}}}};
  assign cxmqpotm = 'bx01;
endmodule: dlcuctbxm

module avawpv
  (output tri0 logic [3:1][1:0] xcp [4:4][3:4], output triand logic [3:3][3:2][3:0] d [2:3][3:1]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xcp = xcp;
  assign d = d;
endmodule: avawpv

module qf
  ( output real vipydimjy
  , input bit [2:1][1:4]  gjpcnhflye
  , input supply1 logic [3:1][0:0][1:3] wvazvlujg [3:3][3:1][0:1][0:2]
  , input tri logic km [2:1]
  , input tri logic [0:0][4:3][2:0] lajfvisi [0:2][0:0][3:4]
  );
  
  
  xor nmrhe(rkh, vipydimjy, vipydimjy);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real vipydimjy -> logic vipydimjy
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real vipydimjy -> logic vipydimjy
  
  not tytbqm(y, vipydimjy);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real vipydimjy -> logic vipydimjy
  
  
  // Single-driven assigns
  assign vipydimjy = gjpcnhflye;
  
  // Multi-driven assigns
  assign wvazvlujg = wvazvlujg;
  assign y = rkh;
  assign rkh = gjpcnhflye;
  assign lajfvisi = lajfvisi;
  assign km = km;
endmodule: qf

module ogguzwzcm
  ();
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ogguzwzcm



// Seed after: 12884744023667183840,5224943229413370507
