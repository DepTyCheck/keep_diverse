// Seed: 12435502455885098234,5224943229413370507

module jtto
  ( output logic [2:4]  tghb
  , output bit [1:3][0:4][4:0]  horeb
  , output logic nlhcdmpg [1:1][0:4]
  , output logic [1:4][4:0][3:2]  qpzav
  , input uwire logic [1:0] k [1:4]
  , input tri1 logic [0:1][1:1][3:4] fbr [4:4]
  );
  
  
  and nocqxwwf(yfcwzo, qpzav, myave);
  // warning: implicit conversion of port connection truncates from 40 to 1 bits
  //   logic [1:4][4:0][3:2]  qpzav -> logic qpzav
  
  
  // Single-driven assigns
  assign tghb = '{'b1001,'b0x,'bx};
  assign horeb = myave;
  
  // Multi-driven assigns
  assign myave = qpzav;
  assign yfcwzo = 'bz0x1;
  assign fbr = fbr;
endmodule: jtto

module rjnq
  ( output int grl [3:4][0:4]
  , output supply1 logic [1:1][4:3][1:4] demhs [1:1]
  , output tri logic iqtpr
  , output supply1 logic pc [4:3][3:3]
  );
  
  
  not ebvpbdc(kbzhpmp, iqtpr);
  
  or shmzyv(iqtpr, kyuei, iqtpr);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign pc = '{'{'b100},'{'b110}};
  assign iqtpr = 'bzzzz1;
  assign demhs = demhs;
  assign kbzhpmp = 'bxz;
endmodule: rjnq



// Seed after: 7537652955198507970,5224943229413370507
