// Seed: 1250704759608574705,5224943229413370507

module bshr
  ( output trireg logic [0:1] ziohjtigf [2:3][0:1][0:4]
  , output logic [4:4][1:3]  odjwbm
  , output reg [1:0][0:0] vh [3:0]
  , input int ftp
  , input tri1 logic dohojtia [3:4][2:4][0:3]
  );
  
  
  not ecwnpu(hmfetumeo, odjwbm);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   logic [4:4][1:3]  odjwbm -> logic odjwbm
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: bshr

module hbxeam
  (input tri logic [2:1][2:1][2:0][2:0] y [4:2][2:3]);
  
  
  not nbwkyfkvv(nhqautpl, nhqautpl);
  
  or yt(nhqautpl, nhqautpl, ulmc);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign nhqautpl = nhqautpl;
  assign ulmc = 'b0110;
  assign y = y;
endmodule: hbxeam



// Seed after: 5966397202017030817,5224943229413370507
