// Seed: 5139529512849536609,5224943229413370507

module hoxmszo
  (output logic kzwbxld);
  
  
  xor cegrupjctd(kzwbxld, hjiss, kzwbxld);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hjiss = hjiss;
endmodule: hoxmszo

module pengzxkzm
  ( output uwire logic [4:2][3:2][1:3][4:3] bgsjfdvtmp [3:4][0:0][3:1][3:4]
  , output realtime rjmx
  , input tri logic [3:1][4:2][3:3][1:1] ubinbcvocp [2:1][4:1][1:2]
  , input bit [4:4][0:0][4:0]  s
  , input triand logic [3:1][0:4] vysh [1:3][0:1][3:1][4:3]
  );
  
  
  nand yhmlyan(rjmx, s, advtyc);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic rjmx -> realtime rjmx
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:0][4:0]  s -> logic s
  
  nand diovqsyfq(oki, rjmx, s);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime rjmx -> logic rjmx
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:0][4:0]  s -> logic s
  
  
  // Single-driven assigns
  assign bgsjfdvtmp = bgsjfdvtmp;
  
  // Multi-driven assigns
  assign advtyc = 'bz11;
  assign vysh = vysh;
  assign oki = rjmx;
  assign ubinbcvocp = ubinbcvocp;
endmodule: pengzxkzm

module ylauzh
  ( output tri1 logic chuexfci [0:1]
  , output logic [0:1][1:3][2:0][1:1]  j
  , input longint srjfadtkvx [0:0]
  , input tri1 logic [0:0][2:4] sz [4:4]
  , input supply0 logic [3:1][1:3][3:1] gvvafbagt [1:2]
  );
  
  
  nand tkksft(sdu, sdu, j);
  // warning: implicit conversion of port connection truncates from 18 to 1 bits
  //   logic [0:1][1:3][2:0][1:1]  j -> logic j
  
  and iovsgocd(fh, kk, hlgsr);
  
  not qstzvf(yrghhnem, kk);
  
  and vwaxpowr(e, a, hlgsr);
  
  
  // Single-driven assigns
  assign j = j;
  
  // Multi-driven assigns
  assign sz = '{'{'{'bzz,'bx111,'bz1}}};
  assign kk = j;
  assign hlgsr = j;
  assign sdu = j;
  assign chuexfci = chuexfci;
endmodule: ylauzh

module zavidlwdnw
  (output realtime vudge, input tri0 logic [4:2][3:0][1:0] mvgzj [4:4], input logic [0:1]  dsvonng);
  
  uwire logic [4:2][3:2][1:3][4:3] vxdp [3:4][0:0][3:1][3:4];
  triand logic [3:1][0:4] kwrdfte [1:3][0:1][3:1][4:3];
  tri logic [3:1][4:2][3:3][1:1] fkplxokht [2:1][4:1][1:2];
  
  xor xihbt(vudge, vudge, vudge);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic vudge -> realtime vudge
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime vudge -> logic vudge
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime vudge -> logic vudge
  
  pengzxkzm ndafiigqfp(.bgsjfdvtmp(vxdp), .rjmx(iycmvefu), .ubinbcvocp(fkplxokht), .s(vudge), .vysh(kwrdfte));
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime rjmx -> wire logic iycmvefu
  //
  // warning: implicit conversion of port connection truncates from 64 to 5 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   realtime vudge -> bit [4:4][0:0][4:0]  s
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign fkplxokht = fkplxokht;
  assign kwrdfte = kwrdfte;
  assign iycmvefu = 'b1zz0;
endmodule: zavidlwdnw



// Seed after: 12148350361508476340,5224943229413370507
