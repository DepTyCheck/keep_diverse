// Seed: 4328217436837865606,5224943229413370507

module jxmql
  ( output bit [1:1][1:1]  piwyaujo
  , output bit [1:4]  vbg
  , output bit [2:1] mynydw [1:4]
  , output logic [3:4][0:2] pvewnwv [2:4]
  , input reg [2:0][4:3]  fdg
  , input logic [2:1]  l
  );
  
  
  not ia(sgw, piwyaujo);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:1][1:1]  piwyaujo -> logic piwyaujo
  
  
  // Single-driven assigns
  assign vbg = '{'b101,'b0,'b1010,'b1};
  
  // Multi-driven assigns
  assign sgw = l;
endmodule: jxmql



// Seed after: 8772000035050567921,5224943229413370507
