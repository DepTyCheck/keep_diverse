// Seed: 16166511167027967125,5224943229413370507

module bzvjul
  ( output logic umnsifa
  , output tri logic [0:3][2:1][3:0][3:1] hgolfsc [4:1][4:3][2:0][0:1]
  , output tri1 logic [3:2][4:3][2:4][2:4] uggf [1:2][1:4][1:3]
  , input logic [0:2][4:0] lcmuwbb [4:1]
  , input logic csbpuyvrie
  , input wor logic [3:1][1:2][3:0] dpruted [2:2][3:3][0:0][4:2]
  );
  
  
  not feer(lwqjraa, hey);
  
  nand bxqpxzg(umnsifa, umnsifa, gkgtoq);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign uggf = uggf;
  assign hgolfsc = hgolfsc;
endmodule: bzvjul



// Seed after: 8101242052950840334,5224943229413370507
