// Seed: 8772000035050567921,5224943229413370507

module w
  ( output bit [1:0][0:3]  avmvdvbe
  , output trireg logic [3:1] vunqatensl [1:1][2:0][0:0]
  , input wand logic [0:2][1:2][1:0][4:1] wermg [2:4][3:4][0:3][2:3]
  );
  
  
  not jae(limwsqmh, avmvdvbe);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:0][0:3]  avmvdvbe -> logic avmvdvbe
  
  not zmrccpyqax(exeimw, avmvdvbe);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:0][0:3]  avmvdvbe -> logic avmvdvbe
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: w



// Seed after: 17851572114395631375,5224943229413370507
