// Seed: 11474204464411577390,5224943229413370507

module ej
  (input logic [1:3][4:3][2:1]  vabqjtfx, input reg [1:2]  trytidj);
  
  
  not fsnwim(q, trytidj);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   reg [1:2]  trytidj -> logic trytidj
  
  not qi(q, trytidj);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   reg [1:2]  trytidj -> logic trytidj
  
  not vmsqmlx(rzlovl, qpprbj);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ej

module bxua
  (input wand logic [1:0] cbesexuywn [2:4][0:4][2:4], input logic [2:1] ikocgcwrp [0:0]);
  
  
  not sc(n, n);
  
  and vsdcrd(n, n, n);
  
  not za(kw, n);
  
  not thuoefmadm(aopd, mblvjfwk);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign n = n;
  assign kw = 'bx0;
  assign mblvjfwk = 'bz1x1;
endmodule: bxua

module gdwwamfzc
  ( output realtime uxl [0:1][4:2]
  , input logic ewvkxlk [4:2][1:0][0:2][1:0]
  , input tri1 logic [1:3][2:4][3:3] g [1:4]
  , input tri1 logic [2:4][1:2] sok [2:1]
  , input reg [4:3][0:4]  o
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign g = '{'{'{'{'bz10z},'{'bxz00x},'{'bzx}},'{'{'bzz0},'{'b0},'{'b00}},'{'{'bx00z0},'{'b0},'{'bxx10z}}},'{'{'{'b0},'{'b1z},'{'bxz01}},'{'{'b0z},'{'b11x},'{'b01}},'{'{'bxxxzx},'{'bxx0z0},'{'b00}}},'{'{'{'bzx},'{'b0},'{'b11z1}},'{'{'b0},'{'b0},'{'b10x}},'{'{'bz},'{'bz},'{'bxzzx0}}},'{'{'{'b0},'{'b0011},'{'b1}},'{'{'bxxz},'{'b1x},'{'b0xzzx}},'{'{'bx},'{'bx0z0},'{'b00zzz}}}};
  assign sok = sok;
endmodule: gdwwamfzc



// Seed after: 16048148996110638788,5224943229413370507
