// Seed: 16249125249849326094,5224943229413370507

module l
  (input wire logic [1:0][3:1] nopepacq [3:0][4:3], input logic [1:3][1:4]  rtotwdir, input real ote [4:0], input reg [1:4] jnciwyi [0:0]);
  
  
  nand j(f, rtotwdir, rtotwdir);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [1:3][1:4]  rtotwdir -> logic rtotwdir
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [1:3][1:4]  rtotwdir -> logic rtotwdir
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign nopepacq = nopepacq;
  assign f = rtotwdir;
endmodule: l

module naq
  ( output trireg logic [4:1][1:1][1:2] x [1:1][1:3]
  , input trireg logic [0:0][0:3][4:1] snzcrwmk [2:0][3:2][4:4]
  , input triand logic [4:1][1:1][1:4][2:1] hbremhk [3:3][1:1]
  , input reg [1:2] dqt [3:0][4:4]
  );
  
  reg [1:4] odoo [0:0];
  real xvyczt [4:0];
  wire logic [1:0][3:1] ejbbs [3:0][4:3];
  
  not teicfpwdjc(pjzqcsj, pjzqcsj);
  
  not ei(pjzqcsj, pjzqcsj);
  
  l qmhbzpnv(.nopepacq(ejbbs), .rtotwdir(pjzqcsj), .ote(xvyczt), .jnciwyi(odoo));
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   wire logic pjzqcsj -> logic [1:3][1:4]  rtotwdir
  
  nand zctzfxpzl(pjzqcsj, glo, pjzqcsj);
  
  
  // Single-driven assigns
  assign xvyczt = '{'bx0x,'b0111,'b10011,'b1z11,'bz1x0};
  assign odoo = odoo;
  
  // Multi-driven assigns
  assign snzcrwmk = snzcrwmk;
endmodule: naq

module pvhkdu
  (output tri1 logic [1:0][4:4] hk [3:2][0:3], output shortreal edxvh, input wire logic [0:0][4:0][1:4] udxcp [0:1][0:3]);
  
  reg [1:4] tmbbailos [0:0];
  real kcalll [4:0];
  wire logic [1:0][3:1] bqsvzpiqg [3:0][4:3];
  
  xor tzykku(bsufvghxpf, edxvh, edxvh);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal edxvh -> logic edxvh
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal edxvh -> logic edxvh
  
  nand nc(zdknvrpr, zdknvrpr, edxvh);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal edxvh -> logic edxvh
  
  l avbs(.nopepacq(bqsvzpiqg), .rtotwdir(edxvh), .ote(kcalll), .jnciwyi(tmbbailos));
  // warning: implicit conversion of port connection truncates from 32 to 12 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal edxvh -> logic [1:3][1:4]  rtotwdir
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hk = hk;
  assign bsufvghxpf = 'bxz;
  assign udxcp = udxcp;
  assign bqsvzpiqg = '{'{'{'{'bx,'b11x,'b1},'{'bzz,'b0z11,'bx1x1}},'{'{'b00z,'bzxxz,'bxzzx},'{'bz,'bz0,'bzz10z}}},'{'{'{'b0,'b0z,'b1xx},'{'bx,'bx,'b1}},'{'{'bx,'bz10,'bzx0z1},'{'b0,'bz,'bz1}}},'{'{'{'b1zzx,'b01xz,'b1xzzx},'{'bx0,'bz,'bx}},'{'{'bz1zzx,'bx0,'bx0z00},'{'b0xzz1,'bz,'bz1x0}}},'{'{'{'bx01,'b0,'bx0x},'{'b1zx11,'bzzz,'b1}},'{'{'b1z,'bx1x1z,'b0z},'{'b00xz,'b0,'b1}}}};
  assign zdknvrpr = bsufvghxpf;
endmodule: pvhkdu



// Seed after: 10771971825523251134,5224943229413370507
