// Seed: 7199167342018908936,5224943229413370507

module ugpdfuawz
  (output reg [0:3][3:2]  urj, input tri logic [1:4][3:0][0:4]  lm, input logic [0:3][2:0]  vjftkf);
  
  
  not zbsp(mq, urj);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [0:3][3:2]  urj -> logic urj
  
  or gd(z, vjftkf, z);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [0:3][2:0]  vjftkf -> logic vjftkf
  
  not y(z, j);
  
  xor qtpkq(lm, urj, urj);
  // warning: implicit conversion of port connection expands from 1 to 80 bits
  //   logic lm -> tri logic [1:4][3:0][0:4]  lm
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [0:3][3:2]  urj -> logic urj
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [0:3][3:2]  urj -> logic urj
  
  
  // Single-driven assigns
  assign urj = '{'{'b10z1,'bzz1},'{'b0z1,'b1},'{'b0000,'bz100z},'{'b0xzz0,'b0}};
  
  // Multi-driven assigns
endmodule: ugpdfuawz

module hya
  ();
  
  
  nand qwnfpnthi(blg, aklg, aklg);
  
  nand omlft(colqrcxzx, aklg, natxwjqd);
  
  ugpdfuawz xuo(.urj(ynm), .lm(tphzlswq), .vjftkf(lpe));
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [0:3][3:2]  urj -> wire logic ynm
  //
  // warning: implicit conversion of port connection expands from 1 to 80 bits
  //   wire logic tphzlswq -> tri logic [1:4][3:0][0:4]  lm
  //
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   wire logic lpe -> logic [0:3][2:0]  vjftkf
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign natxwjqd = natxwjqd;
endmodule: hya

module vqffmxs
  ( output logic bsmb
  , output uwire logic ze [3:1]
  , output logic azy [4:2]
  , output supply1 logic [4:2][1:4][3:4] zxlmdzznn [4:4][4:4]
  , input triand logic [4:4][0:0][4:3][4:3] lesrwpgle [3:1][0:3][1:4][2:3]
  , input tri0 logic [1:4][1:3][0:1][1:3] jkaqoo [3:2][0:1][2:4]
  , input logic [0:2]  htz
  );
  
  
  not ns(oiypr, bsmb);
  
  xor urif(bpruss, htz, bsmb);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   logic [0:2]  htz -> logic htz
  
  not jpkkphekin(bsmb, bsmb);
  
  xor s(eqfhymfb, bsmb, oiypr);
  
  
  // Single-driven assigns
  assign ze = ze;
  assign azy = ze;
  
  // Multi-driven assigns
  assign zxlmdzznn = zxlmdzznn;
  assign eqfhymfb = htz;
  assign jkaqoo = jkaqoo;
  assign oiypr = oiypr;
  assign bpruss = 'bz0;
endmodule: vqffmxs

module yfckfpe
  (output shortreal ruychzkei [1:2][1:4]);
  
  
  nand duwqrk(jwcbwhclcf, f, f);
  
  
  // Single-driven assigns
  assign ruychzkei = ruychzkei;
  
  // Multi-driven assigns
  assign f = f;
  assign jwcbwhclcf = 'b10;
endmodule: yfckfpe



// Seed after: 12515504994790153200,5224943229413370507
