// Seed: 10511653021038236114,5224943229413370507

module ooewc
  ( output realtime cgvmer
  , output reg plwlpf
  , output wor logic [0:0] sjmclrfc [3:3][1:3]
  , input tri logic [2:0] qumduroq [1:4][0:0][1:1][4:2]
  );
  
  
  
  // Single-driven assigns
  assign cgvmer = plwlpf;
  assign plwlpf = 'bx1;
  
  // Multi-driven assigns
endmodule: ooewc

module ndm
  ( output supply0 logic t [4:2]
  , output trior logic [4:3][4:1][3:0] mfguyl [0:2][3:2][1:0][1:2]
  , input reg [4:2][4:3][1:2][0:4]  kdu
  , input logic [3:4] ynljm [4:3]
  , input reg [1:3][3:1][3:1][3:4]  exv
  , input bit [2:2][4:4][3:1][2:0]  fxgmxxj
  );
  
  wor logic [0:0] ti [3:3][1:3];
  tri logic [2:0] crlmcfe [1:4][0:0][1:1][4:2];
  
  not dcrcebiuuw(jawz, kdu);
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   reg [4:2][4:3][1:2][0:4]  kdu -> logic kdu
  
  ooewc zn(.cgvmer(jawz), .plwlpf(jawz), .sjmclrfc(ti), .qumduroq(crlmcfe));
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime cgvmer -> wire logic jawz
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ti = '{'{'{'bz},'{'b00x0},'{'bxzz}}};
endmodule: ndm

module y
  ( output logic fhckxxwuzl [4:0]
  , output trireg logic [4:3][4:2] pzukd [1:4][1:4][1:2]
  , output uwire logic [1:4][2:4][4:0][0:1]  hhthdqwj
  , output bit [1:3][3:1]  prdz
  , input wor logic kzqrxm [4:1][3:1][0:3][2:0]
  , input realtime ptlxg
  );
  
  
  not tjuiqeh(hhthdqwj, hhthdqwj);
  // warning: implicit conversion of port connection expands from 1 to 120 bits
  //   logic hhthdqwj -> uwire logic [1:4][2:4][4:0][0:1]  hhthdqwj
  //
  // warning: implicit conversion of port connection truncates from 120 to 1 bits
  //   uwire logic [1:4][2:4][4:0][0:1]  hhthdqwj -> logic hhthdqwj
  
  not bli(wxlhtur, prdz);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:3][3:1]  prdz -> logic prdz
  
  not cuo(ewgoytvx, ptlxg);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime ptlxg -> logic ptlxg
  
  
  // Single-driven assigns
  assign prdz = '{'{'b1100,'b001,'b1},'{'b11011,'b0,'b01},'{'b01,'b00101,'b0}};
  assign fhckxxwuzl = fhckxxwuzl;
  
  // Multi-driven assigns
  assign pzukd = pzukd;
  assign kzqrxm = kzqrxm;
endmodule: y



// Seed after: 16951114285840472668,5224943229413370507
