// Seed: 2111330656417941348,5224943229413370507

module po
  (output reg [0:4]  ogyio);
  
  
  and vfgwahj(ddvxht, ogyio, duoivvzkjk);
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   reg [0:4]  ogyio -> logic ogyio
  
  nand c(ogyio, uun, ogyio);
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   logic ogyio -> reg [0:4]  ogyio
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   reg [0:4]  ogyio -> logic ogyio
  
  or o(kg, vifahjh, vbmkte);
  
  not ckdmcdx(duoivvzkjk, duoivvzkjk);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign duoivvzkjk = 'b1zz0;
  assign vifahjh = ogyio;
  assign uun = ddvxht;
  assign ddvxht = ogyio;
endmodule: po



// Seed after: 18330800851769687519,5224943229413370507
