// Seed: 2896754593950573947,5224943229413370507

module pdsos
  (input supply0 logic [0:0][2:3] flmlbtzukj [3:3][1:2][2:2], input realtime fr, input supply0 logic [1:4][4:2] rte [4:1]);
  
  
  and epoyfhvcfj(mteusmaii, mteusmaii, mteusmaii);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: pdsos

module gfxshnjvue
  ( output wor logic vsot [3:2]
  , output shortint lwfwfzm
  , input tri1 logic [3:4][1:1][1:1][1:0] o [0:1][3:1][3:1][3:4]
  , input tri0 logic [4:4][3:0][0:3][0:2]  wkgdyeg
  , input bit [0:4][4:2][1:4]  xbtzira
  );
  
  
  
  // Single-driven assigns
  assign lwfwfzm = lwfwfzm;
  
  // Multi-driven assigns
  assign vsot = '{'b0x1x,'bz1x};
  assign wkgdyeg = lwfwfzm;
  assign o = o;
endmodule: gfxshnjvue

module gmmg
  ( output reg [3:1][2:0] e [0:2]
  , output logic [4:2] bwvm [0:3]
  , output logic [1:2][1:1] zmnrw [4:2][1:4]
  , input supply1 logic [1:1][3:0][3:0] gxcke [1:0][2:1]
  );
  
  supply0 logic [1:4][4:2] vwbmebj [4:1];
  supply0 logic [0:0][2:3] c [3:3][1:2][2:2];
  
  pdsos ocd(.flmlbtzukj(c), .fr(evcbtupw), .rte(vwbmebj));
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic evcbtupw -> realtime fr
  
  not xqrwhi(evcbtupw, lhfq);
  
  not znwsjighn(quezryirmc, divy);
  
  or ixzbkwmhi(evcbtupw, cjbyr, quezryirmc);
  
  
  // Single-driven assigns
  assign zmnrw = zmnrw;
  assign bwvm = bwvm;
  assign e = '{'{'{'bx0,'b1x0xx,'b0z0zz},'{'bz11zz,'b00,'bxz},'{'bz1z,'b01xz,'bx}},'{'{'bxx11x,'bx1,'b100z},'{'bzx1,'bz,'b0},'{'bzz10,'bz0,'b11}},'{'{'b0,'b1zx01,'bz},'{'bxz,'bxxzz0,'bx01x},'{'b1,'b0z,'b00z}}};
  
  // Multi-driven assigns
  assign divy = evcbtupw;
  assign evcbtupw = evcbtupw;
  assign c = c;
endmodule: gmmg



// Seed after: 14781989141431543639,5224943229413370507
