// Seed: 8063986785082464560,5224943229413370507

module krsxj
  ( output tri logic [3:3][1:1][3:0][4:2]  p
  , output bit [0:3] ez [1:2][0:3]
  , input reg [2:0][2:3][2:1]  rxycyhgcp
  , input logic [1:4][1:3]  pbidzz
  , input supply0 logic [3:1][2:1][3:0][0:0]  wgdtfxd
  );
  
  
  not zm(p, pbidzz);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic p -> tri logic [3:3][1:1][3:0][4:2]  p
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [1:4][1:3]  pbidzz -> logic pbidzz
  
  or kjbbj(hu, p, pbidzz);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   tri logic [3:3][1:1][3:0][4:2]  p -> logic p
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [1:4][1:3]  pbidzz -> logic pbidzz
  
  
  // Single-driven assigns
  assign ez = ez;
  
  // Multi-driven assigns
  assign p = '{'{'{'{'b1,'b10,'b1zx1},'{'bx,'b1000,'b1zxz},'{'bz11z,'bxxx1z,'b0},'{'bxz,'bzz,'bx0}}}};
endmodule: krsxj

module mivb
  ( output uwire logic [0:3][0:3][4:3] dpngmh [0:1]
  , output real xyvdzuiuu [1:3]
  , output tri logic [0:1][0:2][2:2] qnm [4:1]
  , output wor logic [4:1][4:2][4:2] lbmbibq [3:3][2:1]
  );
  
  
  and ruk(tv, rcewh, bnrixr);
  
  and yfpu(rcewh, rcewh, qeeznpy);
  
  not fkjnbe(rcewh, ni);
  
  
  // Single-driven assigns
  assign dpngmh = '{'{'{'{'bzx11x,'bx00},'{'bz,'b11z1},'{'b1,'bz1zx},'{'bzz,'bx}},'{'{'bxzz0x,'b10xxz},'{'b0xx,'bxx0x},'{'bxxx1,'b0zzzz},'{'bx0111,'b0zz}},'{'{'bzxxzx,'b1},'{'bz0,'b00z0z},'{'bz0xxz,'bx11z},'{'b1x01,'b00}},'{'{'bzx,'bx0zzx},'{'bx0,'b10011},'{'b10,'bz0z1},'{'b0zx,'b1}}},'{'{'{'bz1x,'b00},'{'b1x1,'b01x},'{'bzx,'b101x},'{'bz10,'b1110z}},'{'{'b1z0,'b1z},'{'b00xz,'bx1xz},'{'bx,'bz1x},'{'bx10z,'b0}},'{'{'bz,'bzx0x},'{'bx,'b01x10},'{'bxz0,'b11x10},'{'bz100,'bxx1x}},'{'{'bz,'b0x0z0},'{'b0,'b11},'{'b11,'bz0},'{'b1x0z,'b01x}}}};
  assign xyvdzuiuu = '{'b0xz,'bz,'b0};
  
  // Multi-driven assigns
  assign qeeznpy = 'b01z;
  assign bnrixr = 'b11;
  assign rcewh = tv;
  assign lbmbibq = lbmbibq;
  assign qnm = qnm;
endmodule: mivb

module awv
  ( output real fa
  , output bit yuy
  , output realtime jrhes [3:3]
  , output reg [1:4][0:1][1:2][1:2]  gfes
  , input trireg logic [2:3][4:1][1:0] idg [2:2][3:4][0:0][3:2]
  , input bit [0:3][4:4] l [3:0]
  , input reg [1:2][3:4][1:3]  snluep
  , input wand logic yqajwko [0:0]
  );
  
  bit [0:3] dbntdsuyzq [1:2][0:3];
  
  krsxj abinpx(.p(ricp), .ez(dbntdsuyzq), .rxycyhgcp(gcdl), .pbidzz(gcdl), .wgdtfxd(sy));
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   tri logic [3:3][1:1][3:0][4:2]  p -> wire logic ricp
  //
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   wire logic gcdl -> reg [2:0][2:3][2:1]  rxycyhgcp
  //
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   wire logic gcdl -> logic [1:4][1:3]  pbidzz
  //
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   wire logic sy -> supply0 logic [3:1][2:1][3:0][0:0]  wgdtfxd
  
  xor quwhg(skab, nba, wffieejsgb);
  
  and iqqsondwcs(gfes, yuy, mxrildag);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  //   logic gfes -> reg [1:4][0:1][1:2][1:2]  gfes
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit yuy -> logic yuy
  
  nand rpfvi(kkayccjc, wffieejsgb, jcia);
  
  
  // Single-driven assigns
  assign jrhes = '{'b0111z};
  assign yuy = fa;
  assign fa = 'b001x1;
  
  // Multi-driven assigns
  assign kkayccjc = fa;
  assign nba = 'bzx;
  assign ricp = 'b0x11x;
  assign skab = fa;
  assign gcdl = 'bxxz0z;
endmodule: awv



// Seed after: 4110387113029240658,5224943229413370507
