// Seed: 12862203857658725940,5224943229413370507

module cog
  ( output longint xnjbywhgr [0:1][3:1]
  , output tri1 logic lhqrjpmby
  , output supply1 logic [1:4][1:4][0:4] hpwho [4:0][2:2][0:4][1:3]
  , output bit [0:1]  zkb
  );
  
  
  not wk(qexcwosgrn, zkb);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:1]  zkb -> logic zkb
  
  xor c(lhqrjpmby, qexcwosgrn, qexcwosgrn);
  
  
  // Single-driven assigns
  assign xnjbywhgr = xnjbywhgr;
  assign zkb = lhqrjpmby;
  
  // Multi-driven assigns
  assign qexcwosgrn = zkb;
endmodule: cog

module ttjzlqpig
  ();
  
  supply1 logic [1:4][1:4][0:4] apjgwfb [4:0][2:2][0:4][1:3];
  longint lsxykq [0:1][3:1];
  
  xor egstfdrjtw(he, he, he);
  
  cog ttpcpm(.xnjbywhgr(lsxykq), .lhqrjpmby(he), .hpwho(apjgwfb), .zkb(he));
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:1]  zkb -> wire logic he
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign he = 'b0zx1x;
  assign apjgwfb = apjgwfb;
endmodule: ttjzlqpig

module lfwvsrdjqa
  ( output shortreal kwkmjavbpu
  , input triand logic [0:4][3:1][3:0][2:3] eslnxfze [4:4]
  , input reg [3:1][4:1]  gziovo
  , input shortint mdbf
  );
  
  
  nand ovjec(zyx, wq, kwkmjavbpu);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal kwkmjavbpu -> logic kwkmjavbpu
  
  
  // Single-driven assigns
  assign kwkmjavbpu = zyx;
  
  // Multi-driven assigns
  assign wq = zyx;
  assign eslnxfze = eslnxfze;
  assign zyx = kwkmjavbpu;
endmodule: lfwvsrdjqa

module pcrxa
  ( output supply1 logic zmruo
  , output wor logic [1:2] ptef [1:3][3:2]
  , output tri1 logic [0:0][0:2][0:2] wakkmi [1:0][4:0][4:2]
  , output supply0 logic [4:1][0:3][0:0] ovpiqaizik [4:4]
  , input realtime q [1:1][3:4]
  );
  
  
  and flpmpnqcvo(syfovhglc, zmruo, zmruo);
  
  not obdcqto(k, k);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign zmruo = 'b1z01;
  assign syfovhglc = 'b11x0;
  assign ptef = ptef;
endmodule: pcrxa



// Seed after: 2896754593950573947,5224943229413370507
