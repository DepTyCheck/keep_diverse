// Seed: 13147908407365310562,5224943229413370507

module jpjxlmbd
  (output real vh [0:0], input bit chpnbl, input bit [1:3][2:4]  d, input logic t);
  
  
  
  // Single-driven assigns
  assign vh = '{'b1zzx};
  
  // Multi-driven assigns
endmodule: jpjxlmbd



// Seed after: 2111330656417941348,5224943229413370507
