// Seed: 4710340899852046314,5224943229413370507

module pzqhb
  ( output wand logic [1:1][2:3][4:4][1:4]  tx
  , output wor logic [0:2][4:3] bpvvuer [3:1][1:1][0:4]
  , output bit [0:0][3:1][4:2]  itvf
  , input byte thtrwq
  );
  
  
  not pgklhcvp(tx, tx);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  //   logic tx -> wand logic [1:1][2:3][4:4][1:4]  tx
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   wand logic [1:1][2:3][4:4][1:4]  tx -> logic tx
  
  
  // Single-driven assigns
  assign itvf = '{'{'{'b0,'b11000,'b01},'{'b010,'b0100,'b01},'{'b0110,'b0011,'b10010}}};
  
  // Multi-driven assigns
  assign bpvvuer = bpvvuer;
  assign tx = '{'{'{'{'b011,'bz,'bz11,'bz0}},'{'{'bx1z,'bx0,'b0x,'bz}}}};
endmodule: pzqhb



// Seed after: 17125441217482363648,5224943229413370507
