// Seed: 16048148996110638788,5224943229413370507

module h
  ( output bit [3:2][1:2][4:3][0:2]  hls
  , output wor logic [2:3][0:3][3:3] vnlf [3:3][3:2]
  , input realtime niydfqmzc
  , input bit [2:1][4:4][2:3]  jv
  , input reg [3:4]  chcbwwsd
  );
  
  
  not brkfjelvc(lnwj, niydfqmzc);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime niydfqmzc -> logic niydfqmzc
  
  
  // Single-driven assigns
  assign hls = '{'{'{'{'b0,'b110,'b10110},'{'b0,'b0111,'b1}},'{'{'b00,'b1010,'b1110},'{'b1,'b10011,'b00111}}},'{'{'{'b10111,'b11,'b01010},'{'b0101,'b0,'b011}},'{'{'b10000,'b01010,'b10000},'{'b0,'b111,'b10001}}}};
  
  // Multi-driven assigns
  assign lnwj = 'b11x;
  assign vnlf = vnlf;
endmodule: h

module lahls
  (output reg [2:3]  hpsdhxfwr, output logic f, output tri0 logic [0:2][4:2][3:4]  r, output wor logic [2:0] xio [3:0][2:0][3:3]);
  
  
  not fibi(hpsdhxfwr, kcv);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic hpsdhxfwr -> reg [2:3]  hpsdhxfwr
  
  
  // Single-driven assigns
  assign f = r;
  
  // Multi-driven assigns
  assign r = '{'{'{'bx1,'b110z},'{'b1x00,'bx01},'{'bxx11,'bxxz1x}},'{'{'b0x0z0,'bx1x10},'{'b0xx0,'b01x},'{'bxzxx1,'b1x}},'{'{'b0,'b1},'{'bz1,'b101x},'{'bxxx0,'bx}}};
endmodule: lahls

module jlps
  (output bit tjsyuwsh [3:3], input bit [1:4][2:3][3:1][2:3]  b, input tri0 logic [1:1][0:2] lzvynl [3:1][1:0][1:4]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: jlps



// Seed after: 17479392991164232186,5224943229413370507
