// Seed: 3807221459878586453,5224943229413370507

module edfjhvag
  (output trireg logic [1:0] gcvagey [0:3][4:4]);
  
  
  xor mruvn(j, spdtrsqktq, v);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign v = 'b10;
  assign gcvagey = gcvagey;
endmodule: edfjhvag

module uvyaglpo
  ( output logic [4:4] zg [0:0]
  , input logic yxz [2:0]
  , input triand logic [3:3][1:4] pwfi [1:0][1:2][2:4][1:4]
  , input bit [4:3][3:0] roc [2:3]
  );
  
  trireg logic [1:0] kfevhzqu [0:3][4:4];
  
  xor aajf(iwqtixxsg, iwqtixxsg, iwqtixxsg);
  
  edfjhvag mu(.gcvagey(kfevhzqu));
  
  not uhfjajirr(djnapfjwb, clu);
  
  
  // Single-driven assigns
  assign zg = zg;
  
  // Multi-driven assigns
  assign djnapfjwb = 'bx;
  assign pwfi = pwfi;
endmodule: uvyaglpo

module quzcw
  (output logic [0:4][1:4][2:1] wj [0:0], output reg [3:1][2:4]  cqcsz, input tri1 logic xxqgdprkbc [3:3], input reg [4:4]  epko);
  
  logic [4:4] hxp [0:0];
  bit [4:3][3:0] fb [2:3];
  bit [4:3][3:0] rdfggnn [2:3];
  triand logic [3:3][1:4] zqmngw [1:0][1:2][2:4][1:4];
  logic c [2:0];
  
  uvyaglpo kmhffuz(.zg(hxp), .yxz(c), .pwfi(zqmngw), .roc(rdfggnn));
  
  nand pxkv(cqcsz, epko, cm);
  // warning: implicit conversion of port connection expands from 1 to 9 bits
  //   logic cqcsz -> reg [3:1][2:4]  cqcsz
  
  uvyaglpo bofoivt(.zg(xxqgdprkbc), .yxz(c), .pwfi(zqmngw), .roc(fb));
  
  or rflqlilg(cm, cm, cqcsz);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  //   reg [3:1][2:4]  cqcsz -> logic cqcsz
  
  
  // Single-driven assigns
  assign c = '{'bz01,'b1zx,'bx};
  assign fb = rdfggnn;
  assign rdfggnn = rdfggnn;
  assign wj = wj;
  
  // Multi-driven assigns
  assign zqmngw = zqmngw;
  assign xxqgdprkbc = xxqgdprkbc;
  assign cm = epko;
endmodule: quzcw

module bzoo
  (output bit [4:3][3:0]  nfeep, input logic p, input wire logic [2:2][2:4]  wxhjft, input trireg logic zm [0:4]);
  
  logic [4:4] khxn [0:0];
  trireg logic [1:0] j [0:3][4:4];
  bit [4:3][3:0] zqngtgnc [2:3];
  triand logic [3:3][1:4] quiklp [1:0][1:2][2:4][1:4];
  logic ht [2:0];
  
  edfjhvag k(.gcvagey(j));
  
  uvyaglpo z(.zg(khxn), .yxz(ht), .pwfi(quiklp), .roc(zqngtgnc));
  
  edfjhvag ejvkddl(.gcvagey(j));
  
  or blouf(cqwtxy, nfeep, lapdcvg);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:3][3:0]  nfeep -> logic nfeep
  
  
  // Single-driven assigns
  assign nfeep = nfeep;
  assign ht = '{'bzx00,'bxz1,'b1};
  assign zqngtgnc = '{'{'{'b10,'b1,'b1011,'b10001},'{'b0010,'b01,'b110,'b11010}},'{'{'b0010,'b01,'b10101,'b10},'{'b01,'b1,'b01,'b11110}}};
  
  // Multi-driven assigns
  assign cqwtxy = nfeep;
  assign quiklp = quiklp;
  assign zm = '{'bz0z,'b000,'bz00,'bz1,'bz1x};
endmodule: bzoo



// Seed after: 2626356992014929702,5224943229413370507
