// Seed: 12351719311329769388,5224943229413370507

module stwwpizvtu
  (output reg [3:3][4:3][0:2][3:4]  jf, input bit [3:3][4:4][0:4][4:3]  hwlguuruy, input shortreal kqot [0:3][3:0][3:0]);
  
  
  not ofnwwxfjok(gzvhpp, jf);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [3:3][4:3][0:2][3:4]  jf -> logic jf
  
  
  // Single-driven assigns
  assign jf = '{'{'{'{'bx,'bz101},'{'bz0x,'bx},'{'bz0,'bx}},'{'{'bxz1,'bzz},'{'bxx,'b1},'{'bzxz00,'b10}}}};
  
  // Multi-driven assigns
  assign gzvhpp = hwlguuruy;
endmodule: stwwpizvtu

module winrryyl
  (output triand logic [4:3][4:4] xxhhbq [0:4], input tri0 logic [1:2][1:2]  szh, input reg [2:4]  a);
  
  
  xor dwohodg(szh, szh, szh);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic szh -> tri0 logic [1:2][1:2]  szh
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   tri0 logic [1:2][1:2]  szh -> logic szh
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   tri0 logic [1:2][1:2]  szh -> logic szh
  
  nand mvg(szh, a, xnosopuf);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic szh -> tri0 logic [1:2][1:2]  szh
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   reg [2:4]  a -> logic a
  
  not wmblhmfnoq(szh, dxsyhbveku);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic szh -> tri0 logic [1:2][1:2]  szh
  
  not vc(qntvspx, lm);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xxhhbq = xxhhbq;
endmodule: winrryyl



// Seed after: 3136145052316200612,5224943229413370507
