// Seed: 7162295197203263696,5224943229413370507

module kgxcgigqup
  (output triand logic [3:3][2:4][1:2][3:4] tvduidrmj [4:2][2:0][3:2][1:0], output bit [2:1][4:1][1:3][0:1]  iem, input logic xyr [4:2]);
  
  
  
  // Single-driven assigns
  assign iem = '{'{'{'{'b1000,'b1},'{'b0,'b01000},'{'b10111,'b01}},'{'{'b0,'b0},'{'b0111,'b1},'{'b1110,'b010}},'{'{'b10,'b001},'{'b101,'b0},'{'b1100,'b1111}},'{'{'b10,'b11},'{'b11000,'b00000},'{'b11,'b000}}},'{'{'{'b010,'b110},'{'b00000,'b0},'{'b0111,'b00001}},'{'{'b00,'b110},'{'b000,'b111},'{'b101,'b1011}},'{'{'b0,'b1},'{'b001,'b1011},'{'b000,'b0}},'{'{'b001,'b10},'{'b11111,'b00},'{'b11100,'b1100}}}};
  
  // Multi-driven assigns
  assign tvduidrmj = tvduidrmj;
endmodule: kgxcgigqup

module a
  (output logic [2:0][4:3] xfzettg [4:2][4:3], input reg wmhm [1:4], input tri1 logic [2:2][3:4][2:0] xedghhiksx [2:2]);
  
  
  xor xrmp(afwvhhl, afwvhhl, ipnkxqhuvf);
  
  nand jscqdsde(vpo, afwvhhl, afwvhhl);
  
  
  // Single-driven assigns
  assign xfzettg = '{'{'{'{'b01,'bz},'{'bx000z,'bz},'{'bx10,'b0zxx0}},'{'{'b10,'b11x0},'{'bz1,'b10},'{'bz0z00,'b0xz0}}},'{'{'{'b1zx1x,'b001xz},'{'bx,'bz011x},'{'bx01,'b01zz}},'{'{'b00xz,'bzzz0},'{'bz0xx1,'bz},'{'bzzx0,'b010}}},'{'{'{'b1zzxx,'bxx00x},'{'bzx000,'b1},'{'b1z,'b00zzz}},'{'{'bzx11,'b0zxz},'{'bxx1z,'b1},'{'bxx,'bz}}}};
  
  // Multi-driven assigns
  assign xedghhiksx = '{'{'{'{'bzz11z,'b0,'b0z11},'{'bx0,'bx,'bzz00}}}};
  assign ipnkxqhuvf = ipnkxqhuvf;
  assign afwvhhl = 'b0xx11;
  assign vpo = afwvhhl;
endmodule: a



// Seed after: 153379833403067118,5224943229413370507
