// Seed: 17125441217482363648,5224943229413370507

module mrgua
  (output wire logic thw [3:1][2:1]);
  
  
  and y(ookyqm, ookyqm, vww);
  
  xor dmceol(cdvxmj, adrrhzuqk, ookyqm);
  
  not npsosq(ookyqm, rxrtkfevq);
  
  not uuuicvpr(ookyqm, pbyshxigav);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign thw = thw;
  assign pbyshxigav = ookyqm;
  assign ookyqm = adrrhzuqk;
endmodule: mrgua

module hnpwiuxfs
  (input logic [1:1][4:4][0:0]  dkwhfl, input logic [3:2]  byfhqnzhun, input uwire logic [1:4][2:2][1:3][1:4] vfpr [2:1][4:0][4:2]);
  
  wire logic pcdk [3:1][2:1];
  
  not vy(ilfor, byfhqnzhun);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   logic [3:2]  byfhqnzhun -> logic byfhqnzhun
  
  mrgua odvesjrhn(.thw(pcdk));
  
  xor pflrrmwhb(xdo, xdo, byfhqnzhun);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   logic [3:2]  byfhqnzhun -> logic byfhqnzhun
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ilfor = ilfor;
endmodule: hnpwiuxfs



// Seed after: 17257244788408976843,5224943229413370507
