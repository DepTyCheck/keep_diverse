// Seed: 6917880248887914702,5224943229413370507

module xlageesnhm
  (input supply1 logic [0:3] rbtf [3:1][4:1][0:1][4:0]);
  
  
  not wsnqgdna(mwgu, tiymwvdbz);
  
  xor utwed(tiymwvdbz, jluyrh, tiymwvdbz);
  
  not shae(a, zlnrg);
  
  nand x(mwgu, tiymwvdbz, idsxy);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign mwgu = 'b0xz;
endmodule: xlageesnhm

module sbbgwz
  (output shortint fmq, input reg vehtarrw, input uwire logic [2:2][4:4][4:2][3:4]  sopooy);
  
  
  
  // Single-driven assigns
  assign fmq = fmq;
  
  // Multi-driven assigns
endmodule: sbbgwz

module kuo
  (output reg [3:3][3:0][3:1]  ahf, output supply0 logic [0:3][3:4][4:1][3:2] ferzq [0:2][0:3]);
  
  
  
  // Single-driven assigns
  assign ahf = '{'{'{'bx00z0,'b1z01,'bzz11},'{'b0xx,'bx0,'bzzz1},'{'b1,'b01xx,'b1z011},'{'bz1,'b011,'b1z001}}};
  
  // Multi-driven assigns
  assign ferzq = ferzq;
endmodule: kuo



// Seed after: 17572085871436220380,5224943229413370507
