// Seed: 4242792654842282648,5224943229413370507

module maowwsld
  ( output supply0 logic [1:2][1:2][3:3] jjn [0:1][0:4][0:4][2:3]
  , output supply1 logic [2:3] yhkkoz [4:1][4:4]
  , input longint jid [0:1][3:1]
  , input integer efammlu
  , input reg [4:0][3:4] urzraf [4:4]
  );
  
  
  not k(txxmvkisci, x);
  
  nand igmczvv(heczc, x, heczc);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: maowwsld

module un
  ( output real fnfti [3:0][0:3]
  , output trireg logic [0:3][4:0][2:2] hmzwr [2:2][3:1]
  , output wire logic [2:0][1:3] kfnf [4:2][0:2][2:4][1:4]
  , input wire logic [0:1][0:4][1:3] grnga [1:0][2:1][4:1][3:2]
  );
  
  supply0 logic [1:2][1:2][3:3] vtbu [0:1][0:4][0:4][2:3];
  supply1 logic [2:3] bjbfewjvr [4:1][4:4];
  supply0 logic [1:2][1:2][3:3] xzdafnxlpo [0:1][0:4][0:4][2:3];
  reg [4:0][3:4] h [4:4];
  reg [4:0][3:4] znfsessr [4:4];
  longint uiebrlhvhy [0:1][3:1];
  reg [4:0][3:4] ufg [4:4];
  longint ctu [0:1][3:1];
  
  maowwsld bfuftdgtkp(.jjn(xzdafnxlpo), .yhkkoz(bjbfewjvr), .jid(ctu), .efammlu(tfngp), .urzraf(ufg));
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic tfngp -> integer efammlu
  
  maowwsld oadqisa(.jjn(vtbu), .yhkkoz(bjbfewjvr), .jid(uiebrlhvhy), .efammlu(tfngp), .urzraf(znfsessr));
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic tfngp -> integer efammlu
  
  maowwsld rpn(.jjn(xzdafnxlpo), .yhkkoz(bjbfewjvr), .jid(ctu), .efammlu(tfngp), .urzraf(h));
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic tfngp -> integer efammlu
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: un

module wuegjfhui
  ( output logic wclfvdmztg [2:4][0:2][1:0]
  , output bit [0:0][2:1]  t
  , input tri1 logic [2:0][1:4][2:4][3:0]  ksnqp
  , input trior logic k [1:0][0:3]
  );
  
  wire logic [2:0][1:3] naaruqx [4:2][0:2][2:4][1:4];
  trireg logic [0:3][4:0][2:2] ahkxtshxp [2:2][3:1];
  real hehluyz [3:0][0:3];
  wire logic [0:1][0:4][1:3] lbyd [1:0][2:1][4:1][3:2];
  
  un vnvn(.fnfti(hehluyz), .hmzwr(ahkxtshxp), .kfnf(naaruqx), .grnga(lbyd));
  
  
  // Single-driven assigns
  assign wclfvdmztg = wclfvdmztg;
  assign t = t;
  
  // Multi-driven assigns
  assign ksnqp = t;
  assign k = k;
  assign naaruqx = naaruqx;
  assign lbyd = lbyd;
endmodule: wuegjfhui

module devrpll
  ( output real fjtmw [3:4][1:3][2:3]
  , output logic j [1:2][4:0]
  , output reg hicx
  , output logic [0:2]  wpmtkn
  , input supply1 logic [1:1][2:2][3:3] irooeoyshu [1:1][0:1][0:1]
  , input shortint cvftqt
  );
  
  supply1 logic [2:3] cnnitfwwh [4:1][4:4];
  supply0 logic [1:2][1:2][3:3] pipjsqg [0:1][0:4][0:4][2:3];
  reg [4:0][3:4] m [4:4];
  longint hfr [0:1][3:1];
  
  not crniok(hjtsg, wpmtkn);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   logic [0:2]  wpmtkn -> logic wpmtkn
  
  maowwsld moybawvpx(.jjn(pipjsqg), .yhkkoz(cnnitfwwh), .jid(hfr), .efammlu(cvftqt), .urzraf(m));
  // warning: implicit conversion of port connection expands from 16 to 32 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint cvftqt -> integer efammlu
  
  
  // Single-driven assigns
  assign hicx = 'b10x1;
  assign j = '{'{'b0001x,'bz1,'bx,'b1z1zz,'b0z110},'{'bxxx,'bx0z,'bx1,'bzxx,'bz11}};
  assign fjtmw = '{'{'{'b011z,'bz100z},'{'bx0zz,'bxzz0},'{'bz,'b0x10}},'{'{'bzzz1,'b1xz},'{'b10x1,'b10z},'{'b0101,'bx}}};
  
  // Multi-driven assigns
endmodule: devrpll



// Seed after: 561102826984812543,5224943229413370507
