// Seed: 9771841626331172684,5224943229413370507

module qgp
  (output tri0 logic [4:1][1:4] xb [1:0][4:4][3:3][4:1], output time pj [4:3][0:3][0:4], output int cj [0:1], output shortreal ilifh);
  
  
  nand l(fyoc, a, jssrigheg);
  
  
  // Single-driven assigns
  assign ilifh = 'bxz;
  assign cj = '{'b1001,'b0};
  assign pj = '{'{'{'b1z0,'b1x,'bzzzzx,'bxx0z,'bzz1xx},'{'bxx,'b0,'bxz1x,'bx,'bzx},'{'b1zzxz,'b1z,'bxz00,'b0xx0x,'b11111},'{'bx01x,'b1x101,'b1x,'b1,'b1x1z}},'{'{'b01,'b0,'b10,'bzz1x,'b1xz1x},'{'b1xxxz,'b0,'b0001x,'bxz0z,'bxx},'{'b1xx0x,'bz010,'bxx111,'bx0,'b0},'{'bz0,'bz111,'bz010z,'b00,'bzz}}};
  
  // Multi-driven assigns
  assign fyoc = jssrigheg;
endmodule: qgp

module w
  (output bit [0:1][4:2][3:3]  bgxejzt, output shortint vd [1:2][4:4], input shortint ooyxw);
  
  
  not ajssmucij(bgxejzt, bgxejzt);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic bgxejzt -> bit [0:1][4:2][3:3]  bgxejzt
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:1][4:2][3:3]  bgxejzt -> logic bgxejzt
  
  xor xtjjau(bchqlunyf, bgxejzt, bchqlunyf);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:1][4:2][3:3]  bgxejzt -> logic bgxejzt
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign bchqlunyf = 'b110;
endmodule: w



// Seed after: 8037307645434483667,5224943229413370507
