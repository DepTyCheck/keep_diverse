// Seed: 12884744023667183840,5224943229413370507

module lepsswaod
  ( output trior logic [3:4][3:0][0:4][2:0] vqr [4:1][4:4][3:1][0:2]
  , output bit [2:4][0:1]  p
  , input realtime prhpexde
  , input bit [4:3][3:3][1:1]  dids
  );
  
  
  nand o(p, p, prhpexde);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic p -> bit [2:4][0:1]  p
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][0:1]  p -> logic p
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime prhpexde -> logic prhpexde
  
  not saxipbk(yqrtlr, kssrtwy);
  
  not a(kssrtwy, veq);
  
  and zppl(blhsfjele, prhpexde, p);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime prhpexde -> logic prhpexde
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][0:1]  p -> logic p
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: lepsswaod



// Seed after: 7199167342018908936,5224943229413370507
