// Seed: 11249369895174539472,5224943229413370507

module qixzztrj
  ( output real wshbfy
  , input tri logic i [0:2][4:4][1:0]
  , input logic [2:2]  dlw
  , input supply0 logic [2:1][4:2][3:4] dijl [2:3][3:1]
  );
  
  
  
  // Single-driven assigns
  assign wshbfy = 'b01xx;
  
  // Multi-driven assigns
  assign i = '{'{'{'b10z0,'bx}},'{'{'b0z00,'bz}},'{'{'bxzz,'b1x0x}}};
  assign dijl = dijl;
endmodule: qixzztrj

module sjpwkbtd
  (output trireg logic [4:2][0:0] yn [1:4][3:0][1:3][2:4]);
  
  supply0 logic [2:1][4:2][3:4] cyom [2:3][3:1];
  tri logic rimmzbau [0:2][4:4][1:0];
  
  not yd(o, o);
  
  not go(gtiinfsnz, o);
  
  qixzztrj qzhj(.wshbfy(imxhvgjfue), .i(rimmzbau), .dlw(o), .dijl(cyom));
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real wshbfy -> wire logic imxhvgjfue
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: sjpwkbtd

module sxwgulfyg
  ( output shortreal fnxlubz [4:4][2:4]
  , output tri0 logic [2:1][4:1] sta [1:2][4:4][0:3]
  , output logic [2:2] hobwi [1:2]
  , output supply0 logic [1:0]  todqsmsk
  , input triand logic [3:2][1:1] l [2:2]
  , input tri logic [2:3][3:4][4:2] uhnpnxsan [4:1][4:1][1:3][3:0]
  );
  
  
  
  // Single-driven assigns
  assign fnxlubz = fnxlubz;
  assign hobwi = '{'{'bxz0z0},'{'b1x0z}};
  
  // Multi-driven assigns
  assign uhnpnxsan = uhnpnxsan;
  assign todqsmsk = todqsmsk;
  assign l = l;
endmodule: sxwgulfyg



// Seed after: 1397666190550205442,5224943229413370507
