// Seed: 16778707474574903195,5224943229413370507

module rup
  ( output int htrj [1:3]
  , output shortint ztc [4:4]
  , output logic [1:3][4:3][2:2]  yu
  , output supply1 logic [3:0][4:4][3:4][1:1] ih [1:0][0:3][4:1]
  , input wand logic [3:1][1:1][1:3] ingjwa [0:1][3:1][1:1][0:2]
  , input trireg logic civpygzr [1:2][1:4][0:3][2:2]
  );
  
  
  not rg(npvhtew, yu);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [1:3][4:3][2:2]  yu -> logic yu
  
  not zamfqkiqiw(iimh, yu);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [1:3][4:3][2:2]  yu -> logic yu
  
  not kvankdwi(yu, yu);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   logic yu -> logic [1:3][4:3][2:2]  yu
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [1:3][4:3][2:2]  yu -> logic yu
  
  xor emjdgsmm(iimh, iimh, ptfl);
  
  
  // Single-driven assigns
  assign htrj = htrj;
  assign ztc = ztc;
  
  // Multi-driven assigns
  assign ingjwa = ingjwa;
  assign ptfl = 'b1;
  assign npvhtew = yu;
  assign ih = ih;
endmodule: rup

module etf
  ();
  
  supply1 logic [3:0][4:4][3:4][1:1] rmomocxtgg [1:0][0:3][4:1];
  shortint mlln [4:4];
  int sewpoy [1:3];
  trireg logic hmipco [1:2][1:4][0:3][2:2];
  wand logic [3:1][1:1][1:3] xtaglivh [0:1][3:1][1:1][0:2];
  
  rup tjpwm(.htrj(sewpoy), .ztc(mlln), .yu(isilmybo), .ih(rmomocxtgg), .ingjwa(xtaglivh), .civpygzr(hmipco));
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [1:3][4:3][2:2]  yu -> wire logic isilmybo
  
  nand yke(veu, postiicck, postiicck);
  
  xor troervjfjh(zs, ovgx, vbzjs);
  
  not yztzsnvmak(ovgx, postiicck);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: etf



// Seed after: 10339972513351536850,5224943229413370507
