// Seed: 7537652955198507970,5224943229413370507

module y
  ( output tri logic [3:3][0:4] o [2:0]
  , input uwire logic [1:0][3:3] xyqfvp [1:0][2:4]
  , input byte mnou
  , input logic [1:2] affkruee [3:2][2:0][3:3]
  , input uwire logic [4:3][4:0] kssxdyb [1:2][3:2][3:1]
  );
  
  
  not i(sf, sf);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign o = o;
endmodule: y

module cl
  (output reg [4:0][4:4] uludg [1:4][4:0], output supply0 logic [3:2] tml [1:3]);
  
  
  or jpom(gwhhvcez, gwhhvcez, gwhhvcez);
  
  not jidsrld(ydygjrimfs, gwhhvcez);
  
  not duesnza(gwhhvcez, gwhhvcez);
  
  not ljcwxazp(e, gwhhvcez);
  
  
  // Single-driven assigns
  assign uludg = uludg;
  
  // Multi-driven assigns
  assign ydygjrimfs = 'bx;
  assign gwhhvcez = 'bxx0;
  assign e = 'b1z0;
  assign tml = '{'{'bxzx,'b00},'{'bzxx,'b00zzz},'{'bxz,'bzzx1x}};
endmodule: cl

module akbllfmod
  ( output integer uekinifg
  , output shortint cjk
  , input logic [1:2] mkxmymbtg [0:0][1:1][4:1]
  , input bit [1:2][3:2] jjxk [3:2]
  , input longint bjkmykl
  );
  
  supply0 logic [3:2] ec [1:3];
  reg [4:0][4:4] oiqipl [1:4][4:0];
  
  cl ytud(.uludg(oiqipl), .tml(ec));
  
  nand borclda(fwcru, uekinifg, bjkmykl);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   integer uekinifg -> logic uekinifg
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint bjkmykl -> logic bjkmykl
  
  
  // Single-driven assigns
  assign uekinifg = uekinifg;
  assign cjk = cjk;
  
  // Multi-driven assigns
  assign ec = ec;
  assign fwcru = uekinifg;
endmodule: akbllfmod

module otfcwhzi
  ( output logic [0:4]  juhea
  , output wand logic [3:2][3:4] kwoewliey [1:3]
  , output bit [3:3][4:0][1:2]  gxlesgl
  , output trior logic dthtqh [0:2][4:0][2:0]
  );
  
  
  
  // Single-driven assigns
  assign juhea = juhea;
  assign gxlesgl = juhea;
  
  // Multi-driven assigns
  assign kwoewliey = '{'{'{'bz1xx0,'b01},'{'b0x1,'bxz00}},'{'{'bz,'b011x},'{'b1x1x0,'b01}},'{'{'bx0,'b10x0},'{'bxz0,'b0xz}}};
  assign dthtqh = '{'{'{'b1,'b001z,'b1},'{'b01x11,'b11,'bz0xxz},'{'b01011,'bzz1zx,'b10z},'{'bz10,'b1x1xz,'b0zzz},'{'b0xzz,'bz0,'bx0}},'{'{'bz00,'bx,'bzz0zx},'{'bzxz,'b010,'b1101z},'{'bx0100,'bzx,'b1},'{'bx,'b1z00x,'bzxz11},'{'bxz0xz,'bxzzx,'b01}},'{'{'b11z,'b1x1zz,'bx0111},'{'b1z0zx,'bx11z,'b01},'{'b1zxxz,'b1x00,'b1},'{'bxzzx,'bxxz,'bx1},'{'bz,'bx1,'b01}}};
endmodule: otfcwhzi



// Seed after: 4633840483661197833,5224943229413370507
