// Seed: 17572085871436220380,5224943229413370507

module ycwkot
  (output realtime egt, input real enj, input wire logic [4:1]  uqfbucsj);
  
  
  not kpex(kziyscg, egt);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime egt -> logic egt
  
  or tpufmfav(i, enj, egt);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real enj -> logic enj
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime egt -> logic egt
  
  and wpyyzrg(egt, egt, enj);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic egt -> realtime egt
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime egt -> logic egt
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real enj -> logic enj
  
  or u(uqfbucsj, tnhcu, pbmqu);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic uqfbucsj -> wire logic [4:1]  uqfbucsj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign tnhcu = 'bz0z;
endmodule: ycwkot



// Seed after: 8063986785082464560,5224943229413370507
