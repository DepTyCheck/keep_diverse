// Seed: 12436611882516698977,5224943229413370507

module yicjcnpzyh
  (output bit [1:4][4:0]  o, input uwire logic mdx [2:4], input reg dti);
  
  
  nand udkurid(vgyab, o, bpcadfim);
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][4:0]  o -> logic o
  
  not dnwbmu(hrvegy, vgyab);
  
  not ykdfr(o, o);
  // warning: implicit conversion of port connection expands from 1 to 20 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic o -> bit [1:4][4:0]  o
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][4:0]  o -> logic o
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign bpcadfim = 'b1x;
  assign hrvegy = 'b0z11;
  assign vgyab = 'bzzz;
endmodule: yicjcnpzyh

module qpcocxc
  ( output supply1 logic bmjsudjkj [1:3][1:1][1:3]
  , output reg b [3:2]
  , output supply1 logic [4:3][3:4][0:4] et [4:0][1:3][2:1]
  , input bit ltjnvv
  , input tri1 logic [4:0][3:1] djfpvinesu [0:1]
  );
  
  
  not mxe(ooy, ltjnvv);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit ltjnvv -> logic ltjnvv
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: qpcocxc



// Seed after: 11487342626421313432,5224943229413370507
