// Seed: 5966397202017030817,5224943229413370507

module tn
  (input trior logic [1:4] pztudvrm [1:3][4:1]);
  
  
  not nr(ffzvpjr, natulwhwji);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: tn



// Seed after: 13115324323945111150,5224943229413370507
