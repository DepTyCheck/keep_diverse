// Seed: 13898922656242679089,5224943229413370507

module weseqdrq
  ( output bit y
  , output bit [0:0][4:0]  lpjw
  , input trior logic [2:1] gojirz [2:3][0:3][0:4]
  , input wand logic [0:3] e [4:1][3:0][3:2][3:1]
  , input trior logic [1:3][4:1] hsppoy [3:1][3:0][0:4][4:3]
  );
  
  
  
  // Single-driven assigns
  assign y = 'b001;
  assign lpjw = '{'{'b01,'b1,'b1,'b00111,'b01}};
  
  // Multi-driven assigns
  assign hsppoy = hsppoy;
  assign gojirz = gojirz;
endmodule: weseqdrq



// Seed after: 11791960886729708055,5224943229413370507
