// Seed: 15475924140465045634,5224943229413370507

module cqeevdgtbc
  (output shortreal cuipjjg, output integer qpnrer [2:1], output triand logic [1:0] he [2:1][4:2], input wor logic [0:3] dhxodczmsd [3:4][4:1][1:4]);
  
  
  
  // Single-driven assigns
  assign cuipjjg = cuipjjg;
  assign qpnrer = '{'bzz0z,'b0x};
  
  // Multi-driven assigns
  assign he = '{'{'{'b00xx,'bz},'{'b111z,'b0z0},'{'bx,'bxzxx1}},'{'{'bzz10x,'b11},'{'bz1x11,'bzzx1},'{'b0,'bz10}}};
  assign dhxodczmsd = '{'{'{'{'bxz11z,'b1x,'bz0z01,'bx01x},'{'bx1z,'b1xx0,'bx,'b1},'{'bzz1,'bzxz1,'bzx,'b0x},'{'b0x011,'bz0,'b1,'b1}},'{'{'b1,'b0x11z,'b0z00,'bxx},'{'b1xz0,'b00z00,'b0x00z,'bz0z0},'{'b1x11,'bz1,'bzx11,'b1zzz1},'{'bxx,'bz,'bzx101,'bx1}},'{'{'bx00z0,'bz1zx,'bz0,'b0zxx},'{'bzx,'bz,'b1zz0,'b1x},'{'b11z1,'b1zz,'b0x1,'bx0zz},'{'bzzx0,'b0z,'bxz100,'b0z}},'{'{'bxxzzz,'bxzzx,'b0zz00,'b0xx},'{'bx1,'b00x,'bx0011,'bxx00},'{'b01001,'bxx0,'bz,'b1x0z1},'{'bxx1z,'bxzx,'bx,'bx}}},'{'{'{'b0,'b0z0,'b01zx1,'b10},'{'b0z,'b0,'bx,'b1z},'{'bx011z,'b1z1,'b0xxx,'bx},'{'b0,'b11,'bz0,'b0}},'{'{'bz,'bz1xx1,'bxzzzz,'b11100},'{'b00zzz,'bz0,'b0,'b01},'{'bxzz1,'b0xz,'bxzz0,'b00z},'{'bx1,'bxz,'b1,'bx00}},'{'{'bzz,'bzzxx0,'bxx0,'b01zx1},'{'bx101,'bx1,'b10z,'bz10z1},'{'bxz10z,'b0xx,'bzz10,'bxz1z0},'{'bx,'bx0,'b1,'bxx1x}},'{'{'bx01,'bz0,'b00zz1,'b1},'{'b0x0x1,'bxx0x,'b1xx0z,'b000},'{'bx000z,'b101,'bxz11x,'bxxxz},'{'b1101,'b0x,'bxx,'bx0011}}}};
endmodule: cqeevdgtbc

module weafwu
  ( output logic [1:0][2:0][2:0]  mfvbzefh
  , output bit [1:1] blwbhejl [1:4][2:0]
  , input uwire logic [2:4][4:3][1:4] vzmdcddub [3:1][2:0][3:2]
  , input reg [3:2] zupipp [4:2]
  , input tri1 logic zofvsnfrma [4:3]
  , input tri0 logic [2:3][2:4][1:2][0:4] maqan [0:3][2:0]
  );
  
  integer ep [2:1];
  triand logic [1:0] nipe [2:1][4:2];
  integer yeyoenxnz [2:1];
  wor logic [0:3] oa [3:4][4:1][1:4];
  wor logic [0:3] xbmu [3:4][4:1][1:4];
  
  not etyaomi(mfvbzefh, mfvbzefh);
  // warning: implicit conversion of port connection expands from 1 to 18 bits
  //   logic mfvbzefh -> logic [1:0][2:0][2:0]  mfvbzefh
  //
  // warning: implicit conversion of port connection truncates from 18 to 1 bits
  //   logic [1:0][2:0][2:0]  mfvbzefh -> logic mfvbzefh
  
  cqeevdgtbc axvcpotc(.cuipjjg(cmrxyfqme), .qpnrer(yeyoenxnz), .he(nipe), .dhxodczmsd(xbmu));
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal cuipjjg -> wire logic cmrxyfqme
  
  cqeevdgtbc kawvewamg(.cuipjjg(a), .qpnrer(ep), .he(nipe), .dhxodczmsd(oa));
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal cuipjjg -> wire logic a
  
  or rxhtjavvdn(cmrxyfqme, cmrxyfqme, yczr);
  
  
  // Single-driven assigns
  assign blwbhejl = blwbhejl;
  
  // Multi-driven assigns
  assign cmrxyfqme = mfvbzefh;
  assign xbmu = oa;
endmodule: weafwu

module x
  ( output wor logic stdlj
  , output supply0 logic [0:2][4:2][2:3][3:2] ffjfd [0:3][4:3]
  , output reg [3:4][1:1][3:0][3:2]  lbjxghztub
  , output bit frixpsfv
  , input supply1 logic [4:1][1:3] tqnycxcxu [2:4][1:1][2:4][2:3]
  , input trireg logic [0:4] hmrw [1:0][3:3][0:2][4:0]
  );
  
  
  
  // Single-driven assigns
  assign lbjxghztub = stdlj;
  assign frixpsfv = 'b01;
  
  // Multi-driven assigns
  assign stdlj = lbjxghztub;
  assign tqnycxcxu = tqnycxcxu;
  assign ffjfd = ffjfd;
endmodule: x

module wxcwd
  ( output bit [1:4][3:3][2:4]  gejlcrdml
  , output wire logic [0:1][4:3][0:2][0:4] yddqusmc [0:0][4:3][1:4][0:1]
  , output tri1 logic [3:1]  xe
  , output tri logic eocrrlo [3:0]
  );
  
  
  or lihshiu(gejlcrdml, gejlcrdml, w);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic gejlcrdml -> bit [1:4][3:3][2:4]  gejlcrdml
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][3:3][2:4]  gejlcrdml -> logic gejlcrdml
  
  xor e(dng, gejlcrdml, yqm);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][3:3][2:4]  gejlcrdml -> logic gejlcrdml
  
  and dflk(xe, gejlcrdml, y);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic xe -> tri1 logic [3:1]  xe
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][3:3][2:4]  gejlcrdml -> logic gejlcrdml
  
  or muynxeoodc(dng, gejlcrdml, khnukn);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][3:3][2:4]  gejlcrdml -> logic gejlcrdml
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign eocrrlo = eocrrlo;
  assign w = 'bxxx1;
endmodule: wxcwd



// Seed after: 7475688735560469961,5224943229413370507
