// Seed: 1397666190550205442,5224943229413370507

module cxpwrm
  ( output logic [2:3][0:2][0:4]  fsacb
  , output tri0 logic [3:3][2:4][1:3] ioaihakwgl [4:3][0:1]
  , input realtime tuzwutndbk
  , input bit cch
  , input reg [4:4] e [4:4][2:0][1:2]
  , input logic rbxgsp
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ioaihakwgl = ioaihakwgl;
endmodule: cxpwrm

module cp
  ( output shortint hzmr
  , output reg [1:3][3:2][1:0]  adx
  , output tri logic [4:4][0:1][3:4] dsuxx [3:0][0:4]
  , input tri logic [0:0][0:3]  s
  , input wire logic [1:3][1:0][1:2][2:3] m [0:2]
  );
  
  
  nand gjk(pjoczmeffh, pjghqbc, pjghqbc);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign dsuxx = dsuxx;
  assign pjghqbc = adx;
endmodule: cp

module pgbtxeq
  (output reg [0:1][3:2][1:2] hylnjbin [1:3], output tri1 logic [0:3][4:0][0:3][2:1] ojcaae [1:3], output logic [0:1][0:0]  jop);
  
  
  
  // Single-driven assigns
  assign hylnjbin = '{'{'{'{'b0zx,'b10z},'{'bzz0z,'bz1}},'{'{'b01zz,'bx},'{'bzx,'b1x0}}},'{'{'{'bz0xz,'b0z01},'{'b00x,'bx}},'{'{'b0zxz,'b11zz},'{'bxzz,'bzx}}},'{'{'{'b01,'bx},'{'bxzxx0,'bx}},'{'{'bzzx,'bx0},'{'bx,'bz}}}};
  
  // Multi-driven assigns
  assign ojcaae = ojcaae;
endmodule: pgbtxeq

module i
  (input triand logic [3:4][1:4][4:2][2:3] i [2:1], input tri0 logic [1:3][2:0] hvs [4:2]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign i = i;
  assign hvs = '{'{'{'b0zxz1,'b11x0,'b11xz},'{'b10,'bx01x,'b0x0x},'{'b11x1,'bxzz0x,'b1}},'{'{'b0z0,'b0z,'b0},'{'b110,'b0z,'bx},'{'b1,'b1,'b010z}},'{'{'bx,'b0,'b00x1x},'{'bzx0z,'b0x1z,'b00001},'{'b001,'bz1zz,'b1}}};
endmodule: i



// Seed after: 18015104069983429213,5224943229413370507
