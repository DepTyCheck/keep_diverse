// Seed: 3814454678116103976,5224943229413370507

module kmszxalijl
  (input real ias, input logic [3:2][3:4][2:1][2:4]  fzkhr, input bit uecykthxqm, input logic [2:1][2:1][3:0]  odwwy);
  
  
  and lypuze(xvdmrkj, odwwy, odwwy);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   logic [2:1][2:1][3:0]  odwwy -> logic odwwy
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   logic [2:1][2:1][3:0]  odwwy -> logic odwwy
  
  xor iivrdvkq(iukpcz, odwwy, fzkhr);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   logic [2:1][2:1][3:0]  odwwy -> logic odwwy
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   logic [3:2][3:4][2:1][2:4]  fzkhr -> logic fzkhr
  
  nand ekjtgsp(l, ias, ngwinprm);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real ias -> logic ias
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign l = xvdmrkj;
  assign xvdmrkj = 'b0xx10;
  assign iukpcz = fzkhr;
  assign ngwinprm = odwwy;
endmodule: kmszxalijl

module ksp
  ( output tri1 logic [0:1][4:4][3:3] xi [1:3][0:0][4:2]
  , output bit [3:0][3:2][3:0]  cnffgnt
  , input realtime y
  , input bit [2:1][2:0][0:4][1:1]  tgievctq
  , input longint xfpo [2:0][3:1]
  );
  
  
  not hnlogmw(cnffgnt, cs);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic cnffgnt -> bit [3:0][3:2][3:0]  cnffgnt
  
  not nczlxmc(cs, xxdfeg);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xi = xi;
  assign xxdfeg = 'b110;
  assign cs = 'b010x1;
endmodule: ksp

module kxiqqimkaq
  ( input trireg logic [1:3][3:3] zyn [2:1][1:0]
  , input longint lzapvxnkrx
  , input triand logic [4:1][1:4][3:2] sfjtyjkqrt [2:3][3:0]
  , input trireg logic xivg [3:1][4:1]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign zyn = zyn;
  assign xivg = '{'{'bzz0,'b00z,'bzx,'bx},'{'b00x,'b101,'b011x,'bzz0},'{'bxx1,'b000,'b0,'bx0zx}};
  assign sfjtyjkqrt = sfjtyjkqrt;
endmodule: kxiqqimkaq



// Seed after: 7162295197203263696,5224943229413370507
