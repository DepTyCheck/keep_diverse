// Seed: 14034477015268381597,5224943229413370507

module gfyzlgs
  (input supply1 logic [0:1][1:1] i [1:2][3:2], input wor logic kowj [0:0][1:1]);
  
  
  nand kwtkpvme(wnigpljs, o, lauf);
  
  xor dyyp(o, lauf, lauf);
  
  not irzqgon(f, qet);
  
  or patabty(wnigpljs, wnigpljs, slatr);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: gfyzlgs

module depk
  ( output reg [1:4] voxohtxr [2:4]
  , output shortint vfmydo [4:4]
  , output tri1 logic rnimsfxd [4:1]
  , output triand logic [0:2] grzzgb [2:3][3:1][0:1][3:4]
  , input reg whxc [3:0][0:3]
  );
  
  
  xor cch(hrc, hrc, gzqpufjaj);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rnimsfxd = rnimsfxd;
  assign gzqpufjaj = hrc;
  assign hrc = hrc;
  assign grzzgb = grzzgb;
endmodule: depk



// Seed after: 5433596400001017772,5224943229413370507
