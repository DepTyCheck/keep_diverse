// Seed: 16951114285840472668,5224943229413370507

module lpz
  ( output logic zzwgpiq [2:1][0:0][1:3]
  , output shortreal wgglqwyx
  , output reg [4:3] evzrt [1:2][3:4][3:4]
  , output uwire logic [0:1][3:2]  ehesivlonu
  );
  
  
  or r(gatpdpunj, wgglqwyx, oec);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal wgglqwyx -> logic wgglqwyx
  
  
  // Single-driven assigns
  assign ehesivlonu = wgglqwyx;
  assign zzwgpiq = '{'{'{'b1x110,'bz1,'bx}},'{'{'bx,'bxz,'bxz0x0}}};
  
  // Multi-driven assigns
  assign gatpdpunj = 'b110;
  assign oec = wgglqwyx;
endmodule: lpz

module s
  ( output real yit
  , output longint svjjlzub
  , input supply1 logic [1:2][0:2] oicfqlwsfb [1:0][0:1]
  , input shortreal xug
  , input trior logic [1:0][2:0] buc [2:4][4:4]
  , input uwire logic [0:3][0:3] vwnqivp [0:0]
  );
  
  
  and vethnxmmx(yit, xug, yit);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic yit -> real yit
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal xug -> logic xug
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real yit -> logic yit
  
  
  // Single-driven assigns
  assign svjjlzub = 'b1;
  
  // Multi-driven assigns
  assign oicfqlwsfb = oicfqlwsfb;
  assign buc = '{'{'{'{'bzx1z,'bx,'bzzz},'{'bz,'b0z,'b0}}},'{'{'{'b11,'bzz,'b1x},'{'bxxxz1,'b1,'b000z0}}},'{'{'{'bx1xz,'b00z,'bz1z},'{'b01x,'bx,'b0}}}};
endmodule: s



// Seed after: 3785318144795445061,5224943229413370507
