// Seed: 4633840483661197833,5224943229413370507

module aqlub
  ();
  
  
  xor arhydxg(csbxhanb, izwwqi, izwwqi);
  
  nand twum(jqsme, izwwqi, fru);
  
  not cqc(tfbtq, kucuvqufj);
  
  and wxtwwk(dv, fru, tfbtq);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign izwwqi = 'bxxx0z;
  assign dv = jqsme;
  assign tfbtq = 'b1;
  assign fru = 'b1x0z;
endmodule: aqlub

module u
  (output trior logic [3:2][4:0]  hu);
  
  
  aqlub v();
  
  or ghtiixu(nhypmpjol, hu, cbkcumlrzq);
  // warning: implicit conversion of port connection truncates from 10 to 1 bits
  //   trior logic [3:2][4:0]  hu -> logic hu
  
  or krshllimu(jncos, it, hu);
  // warning: implicit conversion of port connection truncates from 10 to 1 bits
  //   trior logic [3:2][4:0]  hu -> logic hu
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign it = hu;
endmodule: u



// Seed after: 9916430053765975954,5224943229413370507
