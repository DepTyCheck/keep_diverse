// Seed: 9644684484789254430,5224943229413370507

module csayzam
  (output reg [2:2][2:0][3:4][3:4]  ahzwijinq, output supply1 logic [3:0] rseoav [1:2][4:1][2:4], input reg [0:4][3:0][1:3]  ylss);
  
  
  not tyqxzdncc(mgzmjrbx, ylss);
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   reg [0:4][3:0][1:3]  ylss -> logic ylss
  
  
  // Single-driven assigns
  assign ahzwijinq = ahzwijinq;
  
  // Multi-driven assigns
  assign rseoav = rseoav;
  assign mgzmjrbx = 'bz;
endmodule: csayzam



// Seed after: 15853465871684603681,5224943229413370507
