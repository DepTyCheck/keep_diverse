// Seed: 5054388276277724192,5224943229413370507

module w
  (input tri logic kxpuyl, input wire logic [0:0][4:4][1:3] x [2:1][4:1][2:4], input tri logic [4:4] mdbl [1:1][4:4][0:0][2:1]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kxpuyl = 'b1x;
  assign x = x;
endmodule: w

module xppu
  ( output logic [4:4][3:3] fqxpihqrv [3:4][4:3]
  , output shortreal ihsrcdqtcm
  , output tri1 logic [0:4][4:0][0:1][4:0] lsrfnd [3:3]
  , output supply0 logic yknfy [0:4][2:1]
  , input longint xa
  , input supply1 logic [3:4][2:2][1:4] vt [2:3][4:4][1:0]
  );
  
  
  nand fue(ihsrcdqtcm, ihsrcdqtcm, ihsrcdqtcm);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic ihsrcdqtcm -> shortreal ihsrcdqtcm
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal ihsrcdqtcm -> logic ihsrcdqtcm
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal ihsrcdqtcm -> logic ihsrcdqtcm
  
  
  // Single-driven assigns
  assign fqxpihqrv = '{'{'{'{'b1zzx}},'{'{'bxx001}}},'{'{'{'bz}},'{'{'bz}}}};
  
  // Multi-driven assigns
  assign yknfy = '{'{'bxx10,'bx0z},'{'bzx1x,'bzx1},'{'bxxz0,'b01z0},'{'b1011z,'bx},'{'b0x0,'b1}};
  assign lsrfnd = lsrfnd;
  assign vt = vt;
endmodule: xppu

module wnckagub
  (output realtime gn [4:3], output reg jwbcbo, input bit udz, input trireg logic v [4:4][2:3][1:1][1:0]);
  
  
  not pcktu(bbrblfvxex, udz);
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit udz -> logic udz
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign v = v;
  assign bbrblfvxex = jwbcbo;
endmodule: wnckagub

module bm
  ( output trior logic [1:1][2:3][3:2][1:2] ldp [1:2]
  , output logic [1:2][4:4][4:4]  vb
  , output shortreal qqtfyu
  , input wor logic [4:3] tev [0:4][4:3][0:3][4:3]
  , input logic [4:0] rctzvcda [2:4][3:2]
  , input wor logic [0:1][4:4] eumc [4:3][3:2][2:4]
  );
  
  
  
  // Single-driven assigns
  assign qqtfyu = 'b0z1;
  assign vb = vb;
  
  // Multi-driven assigns
  assign tev = tev;
  assign eumc = eumc;
  assign ldp = ldp;
endmodule: bm



// Seed after: 10511653021038236114,5224943229413370507
