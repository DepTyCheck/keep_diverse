// Seed: 9772030656613686378,5224943229413370507

module zbt
  ( output reg [3:3][4:0][4:0]  sppfcx
  , output reg [2:1][2:2] odzcui [2:4][2:3]
  , output reg ih [3:2]
  , input logic [1:4][4:0][2:4][3:3]  hnofwkqokt
  , input shortreal ut
  );
  
  
  xor bomq(ubpjcvid, hnofwkqokt, glbcxw);
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   logic [1:4][4:0][2:4][3:3]  hnofwkqokt -> logic hnofwkqokt
  
  not ueqsm(ihsfhhew, nley);
  
  or q(ubpjcvid, sppfcx, ubpjcvid);
  // warning: implicit conversion of port connection truncates from 25 to 1 bits
  //   reg [3:3][4:0][4:0]  sppfcx -> logic sppfcx
  
  
  // Single-driven assigns
  assign sppfcx = sppfcx;
  
  // Multi-driven assigns
  assign glbcxw = 'b1xxx0;
endmodule: zbt

module t
  ( output wor logic [2:4][3:4][1:0][0:0] nmoovedx [0:1][2:1]
  , output wor logic w [4:3]
  , output longint ptuuvehj
  , input reg qom [0:2]
  , input reg [0:2][3:1] mcxl [2:4]
  );
  
  
  not vnpjbs(hyi, ptuuvehj);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ptuuvehj -> logic ptuuvehj
  
  and jizyj(ptuuvehj, ptuuvehj, ptuuvehj);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic ptuuvehj -> longint ptuuvehj
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ptuuvehj -> logic ptuuvehj
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ptuuvehj -> logic ptuuvehj
  
  not ifielk(aqrxhaxr, ptuuvehj);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ptuuvehj -> logic ptuuvehj
  
  not swtbber(rzhqexd, rzhqexd);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: t

module rjwckj
  (output int axuv, input tri1 logic [1:1]  pkgqotxhu, input reg yxqp);
  
  wor logic xtld [4:3];
  wor logic [2:4][3:4][1:0][0:0] ilczdbmcoj [0:1][2:1];
  reg [0:2][3:1] fads [2:4];
  reg d [0:2];
  
  t bjsu(.nmoovedx(ilczdbmcoj), .w(xtld), .ptuuvehj(qy), .qom(d), .mcxl(fads));
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   longint ptuuvehj -> wire logic qy
  
  nand jms(fugye, axuv, axuv);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int axuv -> logic axuv
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int axuv -> logic axuv
  
  
  // Single-driven assigns
  assign axuv = 'b1;
  assign fads = '{'{'{'bzxzxx,'b0,'b1xx},'{'bzz,'b1zz,'bx1xx},'{'b001xz,'bzz0z,'bxx}},'{'{'b000,'b1x,'b1},'{'b0,'bxx,'b1z000},'{'b101xx,'bx1,'b0}},'{'{'bz0,'b1,'b00zz},'{'b0z,'bx10,'bz1},'{'b0,'b1x1,'bxx}}};
  assign d = d;
  
  // Multi-driven assigns
  assign fugye = 'b0xx1;
  assign xtld = '{'bx,'b11xz};
  assign ilczdbmcoj = ilczdbmcoj;
  assign qy = yxqp;
  assign pkgqotxhu = axuv;
endmodule: rjwckj

module j
  (output logic ya [3:0], input tri0 logic [2:2]  xrwvb);
  
  
  not rnlyedd(xrwvb, xrwvb);
  
  rjwckj vjbsvvsg(.axuv(xrwvb), .pkgqotxhu(xrwvb), .yxqp(cyogzkcnqn));
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int axuv -> tri0 logic [2:2]  xrwvb
  
  
  // Single-driven assigns
  assign ya = '{'b0xzx,'bx1,'bz,'bx};
  
  // Multi-driven assigns
  assign xrwvb = xrwvb;
  assign cyogzkcnqn = 'b0x1x;
endmodule: j



// Seed after: 14034477015268381597,5224943229413370507
