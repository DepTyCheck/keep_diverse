// Seed: 11054676645773098073,5224943229413370507

module f
  ( output logic [2:0][1:2][4:0]  j
  , output real mkxmzauc
  , output wire logic [0:0][1:0][2:4][4:2]  awfh
  , output triand logic wvuaufjsu [0:2][1:2][2:2][4:2]
  , input wand logic [1:3][0:0][0:3][3:2] gsnsst [3:2]
  , input logic [4:3][1:0][0:2][3:3]  grfgwukvia
  );
  
  
  not g(hifi, j);
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  //   logic [2:0][1:2][4:0]  j -> logic j
  
  not o(j, j);
  // warning: implicit conversion of port connection expands from 1 to 30 bits
  //   logic j -> logic [2:0][1:2][4:0]  j
  //
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  //   logic [2:0][1:2][4:0]  j -> logic j
  
  and m(kp, mkxmzauc, j);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real mkxmzauc -> logic mkxmzauc
  //
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  //   logic [2:0][1:2][4:0]  j -> logic j
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign gsnsst = gsnsst;
  assign hifi = 'bz1;
  assign awfh = '{'{'{'{'b0,'b100x,'b0},'{'b0z0,'bx,'bx1zz1},'{'b00,'bz00xz,'b0xzz}},'{'{'bx0z0z,'b0z11x,'bz0x},'{'bx1,'bzz10,'bzx11z},'{'b0,'b0zx01,'b1x1zz}}}};
  assign kp = hifi;
  assign wvuaufjsu = '{'{'{'{'b0,'b101,'bzxz}},'{'{'b0z1z,'bxz,'bx1z}}},'{'{'{'b01zz0,'b1x,'bxxz11}},'{'{'b1xxzz,'b11,'b0x1}}},'{'{'{'b1x0,'bxx1z0,'b00z}},'{'{'bxz01,'b1zxx0,'bz1}}}};
endmodule: f

module vuytqudl
  (output logic tjdos, input shortreal so, input logic [3:3]  sqlgres);
  
  triand logic gmimtojfb [0:2][1:2][2:2][4:2];
  wand logic [1:3][0:0][0:3][3:2] zuk [3:2];
  
  or ayjgqhwkl(dtoxizummi, tjdos, tjdos);
  
  f aip(.j(gplezffgfi), .mkxmzauc(mit), .awfh(qpsaik), .wvuaufjsu(gmimtojfb), .gsnsst(zuk), .grfgwukvia(sqlgres));
  // warning: implicit conversion of port connection truncates from 30 to 1 bits
  //   logic [2:0][1:2][4:0]  j -> wire logic gplezffgfi
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real mkxmzauc -> wire logic mit
  //
  // warning: implicit conversion of port connection truncates from 18 to 1 bits
  //   wire logic [0:0][1:0][2:4][4:2]  awfh -> wire logic qpsaik
  //
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic [3:3]  sqlgres -> logic [4:3][1:0][0:2][3:3]  grfgwukvia
  
  not qozwuofq(duwbnd, so);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal so -> logic so
  
  
  // Single-driven assigns
  assign tjdos = tjdos;
  
  // Multi-driven assigns
  assign dtoxizummi = 'b0x;
endmodule: vuytqudl

module bjlxokj
  (output wire logic [0:0][1:2][4:0]  mzq, output bit [2:1][4:1][3:0]  jvd);
  
  
  not rbkb(mzq, mzq);
  // warning: implicit conversion of port connection expands from 1 to 10 bits
  //   logic mzq -> wire logic [0:0][1:2][4:0]  mzq
  //
  // warning: implicit conversion of port connection truncates from 10 to 1 bits
  //   wire logic [0:0][1:2][4:0]  mzq -> logic mzq
  
  nand xtniqocfzw(mzq, rtlzg, jmlxvqf);
  // warning: implicit conversion of port connection expands from 1 to 10 bits
  //   logic mzq -> wire logic [0:0][1:2][4:0]  mzq
  
  
  // Single-driven assigns
  assign jvd = '{'{'{'b1100,'b10,'b00,'b0},'{'b111,'b0101,'b0,'b010},'{'b111,'b100,'b1,'b00001},'{'b1111,'b0,'b11,'b1}},'{'{'b001,'b010,'b00,'b010},'{'b0,'b10101,'b1101,'b10},'{'b0011,'b11,'b0011,'b1},'{'b01,'b0,'b0,'b010}}};
  
  // Multi-driven assigns
  assign mzq = jmlxvqf;
  assign jmlxvqf = jmlxvqf;
endmodule: bjlxokj

module pxgui
  ( output trireg logic [3:3][0:2] trdywkiduk [1:2]
  , output logic mfa
  , output wand logic owrqvk [2:1][0:2]
  , input supply0 logic [0:1][4:1][1:0] lxpdrhel [3:2][2:2][1:2]
  , input uwire logic szjtvotdfd [0:2][1:4]
  );
  
  
  nand eetzgzdjbd(mfa, sdzqghssnj, n);
  
  bjlxokj l(.mzq(dpnkewi), .jvd(nibxzddc));
  // warning: implicit conversion of port connection truncates from 10 to 1 bits
  //   wire logic [0:0][1:2][4:0]  mzq -> wire logic dpnkewi
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:1][4:1][3:0]  jvd -> wire logic nibxzddc
  
  xor zvtae(fw, pahqpquic, mfa);
  
  nand gfgeczgryi(djhzoqitb, fvjmtl, djhzoqitb);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign trdywkiduk = '{'{'{'b1,'b1zz,'b1}},'{'{'bz0,'b0x1,'bx}}};
  assign dpnkewi = 'b0xxxx;
endmodule: pxgui



// Seed after: 10640103557006565659,5224943229413370507
