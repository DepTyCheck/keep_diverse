// Seed: 11487342626421313432,5224943229413370507

module nvsszjj
  (output reg [1:3][3:2] myvxbpjt [2:3][0:0], output reg [0:4][4:1][2:2]  vlvpz);
  
  
  
  // Single-driven assigns
  assign vlvpz = '{'{'{'b1x1z1},'{'b0z},'{'b1},'{'b0zx00}},'{'{'b110},'{'bz1x0},'{'bx},'{'bx01xx}},'{'{'bx},'{'bzx0zz},'{'b10},'{'bz0xzx}},'{'{'b0},'{'bxx11},'{'b0},'{'bxx1z}},'{'{'bz00},'{'b110},'{'b101x},'{'bzx11x}}};
  
  // Multi-driven assigns
endmodule: nvsszjj



// Seed after: 16910038469795232155,5224943229413370507
