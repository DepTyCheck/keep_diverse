// Seed: 2901206930565052048,5224943229413370507

module qbeilo
  (output reg [0:0][3:0]  vtbmc, output logic [2:0]  cieheyywd, output logic [1:4][3:0]  to);
  
  
  and nkwez(bsqxktxlb, mgczlsp, tjms);
  
  not mlwl(mgczlsp, vtbmc);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   reg [0:0][3:0]  vtbmc -> logic vtbmc
  
  not ghgw(vtbmc, tjms);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic vtbmc -> reg [0:0][3:0]  vtbmc
  
  
  // Single-driven assigns
  assign to = mgczlsp;
  
  // Multi-driven assigns
  assign mgczlsp = tjms;
  assign tjms = 'bz1;
endmodule: qbeilo

module pk
  ( input supply0 logic [1:2][0:2]  ljwyqq
  , input bit [3:0][1:2][4:3][0:4]  uq
  , input trireg logic [4:2][2:0][1:3][0:1] owhzh [0:3]
  , input tri logic roeygk [1:3]
  );
  
  
  nand fekkztnf(bu, ilpnqsc, ilpnqsc);
  
  not yuwpi(pcapqiyvvo, ljwyqq);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   supply0 logic [1:2][0:2]  ljwyqq -> logic ljwyqq
  
  not wfigjuvjwj(ugnng, eltrrh);
  
  not urfves(ugbkx, lfipgbpzuf);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign bu = eltrrh;
  assign owhzh = owhzh;
  assign lfipgbpzuf = 'b1z00x;
  assign ilpnqsc = 'b0x1xx;
  assign pcapqiyvvo = ljwyqq;
endmodule: pk



// Seed after: 10835398777294435853,5224943229413370507
