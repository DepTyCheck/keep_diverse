// Seed: 17479392991164232186,5224943229413370507

module guwjzrog
  (output uwire logic [2:3][2:3]  lbzkcmjz);
  
  
  not nyo(zsgwyptvxd, lbzkcmjz);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   uwire logic [2:3][2:3]  lbzkcmjz -> logic lbzkcmjz
  
  not ocfypyvcj(lbzkcmjz, zsgwyptvxd);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic lbzkcmjz -> uwire logic [2:3][2:3]  lbzkcmjz
  
  xor fnwcleep(zsgwyptvxd, lbzkcmjz, lbzkcmjz);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   uwire logic [2:3][2:3]  lbzkcmjz -> logic lbzkcmjz
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   uwire logic [2:3][2:3]  lbzkcmjz -> logic lbzkcmjz
  
  not fbvbpwmw(zsgwyptvxd, ysimyi);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign zsgwyptvxd = lbzkcmjz;
  assign ysimyi = ysimyi;
endmodule: guwjzrog

module yyw
  (output triand logic fgm [4:2][1:3][4:1], output integer bcyfkxxkjw [0:3], input tri0 logic [2:3]  skfsghq);
  
  
  xor xiec(skfsghq, skfsghq, s);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  //   logic skfsghq -> tri0 logic [2:3]  skfsghq
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri0 logic [2:3]  skfsghq -> logic skfsghq
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: yyw

module uhjurmihkk
  (output realtime f, output int ki, output tri logic [1:0][2:0][3:0] ihlih [0:1], output reg ga [1:4]);
  
  
  
  // Single-driven assigns
  assign f = 'bx0z0;
  
  // Multi-driven assigns
endmodule: uhjurmihkk

module xokp
  ( output tri1 logic [3:1][0:4][2:4] rpsqoq [2:2][3:0][4:0][3:2]
  , output tri logic [2:4][3:0] jmzly [0:3][0:0]
  , output reg [4:1][2:2][0:4]  newrbsy
  , input wand logic [2:4] n [2:3][4:3]
  , input logic [3:2][3:4][1:4][0:4]  ulkvgl
  , input shortreal stvxj
  );
  
  integer qefav [0:3];
  triand logic minmsox [4:2][1:3][4:1];
  reg otja [1:4];
  tri logic [1:0][2:0][3:0] menba [0:1];
  
  uhjurmihkk g(.f(efpayzmmuy), .ki(mocvoy), .ihlih(menba), .ga(otja));
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime f -> wire logic efpayzmmuy
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int ki -> wire logic mocvoy
  
  yyw hnajmther(.fgm(minmsox), .bcyfkxxkjw(qefav), .skfsghq(ulkvgl));
  // warning: implicit conversion of port connection truncates from 80 to 2 bits
  //   logic [3:2][3:4][1:4][0:4]  ulkvgl -> tri0 logic [2:3]  skfsghq
  
  or ih(newrbsy, newrbsy, newrbsy);
  // warning: implicit conversion of port connection expands from 1 to 20 bits
  //   logic newrbsy -> reg [4:1][2:2][0:4]  newrbsy
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   reg [4:1][2:2][0:4]  newrbsy -> logic newrbsy
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   reg [4:1][2:2][0:4]  newrbsy -> logic newrbsy
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: xokp



// Seed after: 8957594518452836278,5224943229413370507
