// Seed: 16910038469795232155,5224943229413370507

module blb
  (output bit [3:4][3:2]  vqzseo, input longint rtbwjrs [0:4][0:2][3:4], input triand logic [4:0][4:3] xac [3:3]);
  
  
  not tnjxloan(vqzseo, vqzseo);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic vqzseo -> bit [3:4][3:2]  vqzseo
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:4][3:2]  vqzseo -> logic vqzseo
  
  not vp(bzij, vi);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign vi = 'b00zz0;
  assign bzij = bzij;
  assign xac = xac;
endmodule: blb

module j
  (input bit f, input reg [0:2]  qel, input bit [4:4][3:2]  ywakf, input shortint eobburb [2:1][0:3]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: j

module pmelh
  (output wire logic [2:3][1:1] lvoiu [4:3], input bit [2:3]  wexmhnj, input reg [1:3][1:4]  wq);
  
  shortint pe [2:1][0:3];
  
  j fygiivtt(.f(wexmhnj), .qel(wexmhnj), .ywakf(o), .eobburb(pe));
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   bit [2:3]  wexmhnj -> bit f
  //
  // warning: implicit conversion of port connection expands from 2 to 3 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3]  wexmhnj -> reg [0:2]  qel
  //
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic o -> bit [4:4][3:2]  ywakf
  
  not ezoilmbz(ffakoxird, wexmhnj);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3]  wexmhnj -> logic wexmhnj
  
  
  // Single-driven assigns
  assign pe = '{'{'b11,'b1100,'b1010,'b11},'{'b0010,'b10,'b10101,'b0}};
  
  // Multi-driven assigns
  assign lvoiu = lvoiu;
  assign o = wexmhnj;
  assign ffakoxird = o;
endmodule: pmelh

module gi
  (input triand logic [1:1][0:0][3:4][2:2]  sm, input shortint ox, input wor logic [2:4][0:4][4:2][1:2] mfjuihupcu [1:3]);
  
  
  not yzxhvtl(h, yilgli);
  
  and w(yilgli, yilgli, h);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign yilgli = 'bx;
  assign sm = '{'{'{'{'bxxzx},'{'bz}}}};
endmodule: gi



// Seed after: 11869620239679120121,5224943229413370507
