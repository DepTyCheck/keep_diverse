// Seed: 8957594518452836278,5224943229413370507

module gujzwjbfin
  (output reg [4:3][4:4][4:1] zcpcmyl [0:2], output shortreal icttocr [0:1]);
  
  
  not ry(eoik, uesiatpbys);
  
  and qimma(zazu, q, j);
  
  nand fkqkxsdkuu(diiichkpi, xufbyw, xufbyw);
  
  or rmd(ow, uesiatpbys, jhragchv);
  
  
  // Single-driven assigns
  assign zcpcmyl = '{'{'{'{'b1zx,'bzx0,'b1zx1,'b10}},'{'{'b01z,'bz1,'b0x,'bzxx00}}},'{'{'{'b111,'b0,'b1z1x0,'b1}},'{'{'b1101z,'b10,'bz1z,'bz0xx0}}},'{'{'{'b0,'b1xz,'b001,'b00}},'{'{'bx1,'bx,'bz0z,'bz}}}};
  assign icttocr = '{'b0x,'bxx00x};
  
  // Multi-driven assigns
  assign diiichkpi = 'b1x0;
  assign zazu = 'b1x0;
endmodule: gujzwjbfin

module mqqweoml
  ( input trireg logic [0:1][0:0] lywrt [3:0][0:4]
  , input uwire logic [3:0][4:1][1:1] pit [1:4][2:0][1:1]
  , input tri logic vdlryzkdp [0:2]
  , input bit [3:1][0:4][2:4] bex [4:3]
  );
  
  
  xor aler(ngznhzcet, x, x);
  
  or oxhzc(ngznhzcet, x, x);
  
  not zwcnshl(x, ngznhzcet);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign x = x;
  assign ngznhzcet = x;
  assign lywrt = '{'{'{'{'bz11},'{'b10xz0}},'{'{'bx0},'{'bx}},'{'{'b1x1zz},'{'b0}},'{'{'bzx0},'{'b1}},'{'{'b100xx},'{'bx}}},'{'{'{'b0xx},'{'b0xx}},'{'{'bx0zz},'{'bzxzx}},'{'{'bz0x},'{'bz}},'{'{'bzxz00},'{'b0z0}},'{'{'b0zx},'{'b111}}},'{'{'{'bxzz},'{'b010}},'{'{'b00z},'{'b101}},'{'{'bx},'{'b1}},'{'{'bxx01z},'{'bxxz0}},'{'{'bx10},'{'b0}}},'{'{'{'bxx001},'{'bxx0}},'{'{'bxxzzx},'{'bx}},'{'{'b1x},'{'b11z10}},'{'{'bxzz1},'{'bxx}},'{'{'bz1zz0},'{'bx}}}};
endmodule: mqqweoml



// Seed after: 16058725124331033669,5224943229413370507
