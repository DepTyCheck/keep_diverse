// Seed: 153379833403067118,5224943229413370507

module lwdzfknhls
  ( output reg [2:3] szwgjbw [0:0][4:0]
  , output bit [1:4][3:3] zqxtwfcllb [0:0][3:4]
  , output triand logic [1:1][2:4][1:3][2:4]  ey
  , output tri1 logic [0:4]  yradqvmqrs
  );
  
  
  not jcvpajdmv(vxnhpcelq, xisopjvqq);
  
  not aewgntbqy(vxnhpcelq, vl);
  
  
  // Single-driven assigns
  assign szwgjbw = szwgjbw;
  assign zqxtwfcllb = '{'{'{'{'b0},'{'b00},'{'b10},'{'b0}},'{'{'b10},'{'b110},'{'b10011},'{'b11}}}};
  
  // Multi-driven assigns
  assign ey = xisopjvqq;
  assign vxnhpcelq = 'bzzx;
  assign yradqvmqrs = ey;
endmodule: lwdzfknhls

module ueuqc
  ( output reg [0:4][1:4][3:0][2:4]  qkjeuz
  , output wire logic [0:0][3:2][4:0] dwkwuhlqup [3:1][0:4][3:3][0:1]
  , output wand logic [3:1][1:2][2:1][2:1] fxzqkrxq [1:4][4:4]
  , output shortreal tbvb
  , input real tc [1:0]
  , input integer vylan [1:3]
  );
  
  
  
  // Single-driven assigns
  assign tbvb = qkjeuz;
  
  // Multi-driven assigns
  assign dwkwuhlqup = dwkwuhlqup;
  assign fxzqkrxq = fxzqkrxq;
endmodule: ueuqc

module koie
  (output supply1 logic zslfxjwymp [2:2][3:3][3:3][0:0], input int gczo [1:0][2:2]);
  
  
  xor jjzduhelrh(ha, ha, wfinmkk);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign zslfxjwymp = zslfxjwymp;
endmodule: koie

module no
  ( output logic [0:0][1:4][3:0] vk [4:1]
  , input wand logic [0:3][3:2][2:4][1:2] qxhjmxyr [0:2][4:2][4:3]
  , input longint bujrjzn [4:1]
  , input wor logic [2:1][2:3] alg [4:4][2:4]
  , input wor logic [0:4] w [4:1][4:3][3:2]
  );
  
  bit [1:4][3:3] lmdjqe [0:0][3:4];
  reg [2:3] hfkzhs [0:0][4:0];
  bit [1:4][3:3] s [0:0][3:4];
  reg [2:3] t [0:0][4:0];
  
  lwdzfknhls rrmmf(.szwgjbw(t), .zqxtwfcllb(s), .ey(egyod), .yradqvmqrs(aminqtrbfs));
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  //   triand logic [1:1][2:4][1:3][2:4]  ey -> wire logic egyod
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   tri1 logic [0:4]  yradqvmqrs -> wire logic aminqtrbfs
  
  lwdzfknhls fiz(.szwgjbw(hfkzhs), .zqxtwfcllb(lmdjqe), .ey(ixgfuhnp), .yradqvmqrs(egyod));
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  //   triand logic [1:1][2:4][1:3][2:4]  ey -> wire logic ixgfuhnp
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   tri1 logic [0:4]  yradqvmqrs -> wire logic egyod
  
  or mv(jdaycjf, egyod, egyod);
  
  
  // Single-driven assigns
  assign vk = vk;
  
  // Multi-driven assigns
  assign egyod = 'bzzxxx;
endmodule: no



// Seed after: 4242792654842282648,5224943229413370507
