// Seed: 10835398777294435853,5224943229413370507

module xlsxtrod
  (output logic oybuzskv [3:0][3:3][4:2], output realtime axjjkk, input trireg logic [4:2][3:4][1:2] dukswtkce [4:0]);
  
  
  and cnpcdindy(axjjkk, axjjkk, axjjkk);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic axjjkk -> realtime axjjkk
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime axjjkk -> logic axjjkk
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime axjjkk -> logic axjjkk
  
  
  // Single-driven assigns
  assign oybuzskv = '{'{'{'bx10x,'bzz,'bx0x}},'{'{'b00,'b0x01,'b1}},'{'{'bx11,'b0zxx1,'b0z}},'{'{'b1x,'bxxz1x,'bx}}};
  
  // Multi-driven assigns
endmodule: xlsxtrod

module vruph
  (input tri logic eqjtgp, input trireg logic [4:2][4:0][1:0]  ztdhnzznd, input logic [2:2]  zqgy, input reg qlekedoe [3:4]);
  
  logic vwtshjh [3:0][3:3][4:2];
  trireg logic [4:2][3:4][1:2] x [4:0];
  
  not puvxcnmxip(hydszzmjao, nfosttrip);
  
  not uqucq(hydszzmjao, nfosttrip);
  
  xlsxtrod pxrgqqixpx(.oybuzskv(vwtshjh), .axjjkk(jctnlndj), .dukswtkce(x));
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime axjjkk -> wire logic jctnlndj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hydszzmjao = 'b1001;
  assign x = x;
  assign nfosttrip = nfosttrip;
  assign ztdhnzznd = nfosttrip;
endmodule: vruph

module tdfd
  (output tri logic [1:3][2:2][2:4] khfbafl [4:3], input realtime qbhy [2:4], input bit [2:1][2:0][2:1][1:3]  jvpxmcglf);
  
  
  or oycllk(fdjctr, fdjctr, fdjctr);
  
  and pggmbz(fdjctr, jvpxmcglf, whe);
  // warning: implicit conversion of port connection truncates from 36 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:1][2:0][2:1][1:3]  jvpxmcglf -> logic jvpxmcglf
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign khfbafl = khfbafl;
  assign whe = 'b110z1;
  assign fdjctr = 'b111;
endmodule: tdfd



// Seed after: 9644684484789254430,5224943229413370507
