// Seed: 10339972513351536850,5224943229413370507

module dojp
  (output logic [0:1][3:4][4:0][1:0]  uhgnn, input bit [4:3]  vzqapi, input bit zlr, input trior logic [2:3][0:3][1:2][0:0]  sepsf);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign sepsf = '{'{'{'{'b0zx},'{'b10xx}},'{'{'b0},'{'bx1x1}},'{'{'b0x011},'{'bz}},'{'{'b010},'{'bz0}}},'{'{'{'bxz},'{'b010}},'{'{'bxzz},'{'bx00}},'{'{'b1zxz0},'{'bz0zxz}},'{'{'bxx0},'{'bz1z1z}}}};
endmodule: dojp



// Seed after: 12034918165399613485,5224943229413370507
