// Seed: 6347729663862269036,5224943229413370507

module ptwxgn
  ( output trior logic [2:4]  r
  , output bit qpzmph [2:1]
  , output bit [0:3][0:1][0:1][4:4]  bvuzha
  , input reg twflb
  , input time per
  , input logic [3:4][1:3]  mk
  , input trior logic [0:2][2:4]  fpkakib
  );
  
  
  or mamdui(mw, r, per);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   trior logic [2:4]  r -> logic r
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  //   time per -> logic per
  
  not xwii(r, r);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic r -> trior logic [2:4]  r
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   trior logic [2:4]  r -> logic r
  
  not wz(r, ahtmj);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic r -> trior logic [2:4]  r
  
  nand ohnpmt(jf, ehtwsaw, zith);
  
  
  // Single-driven assigns
  assign qpzmph = '{'b01001,'b1};
  assign bvuzha = r;
  
  // Multi-driven assigns
  assign mw = r;
  assign ahtmj = 'bzz01;
  assign r = r;
  assign zith = 'b11;
endmodule: ptwxgn

module oqexmpwta
  ( output supply1 logic oxexivok
  , output trireg logic [3:3][3:0]  iurbtodez
  , output wire logic [3:2] in [4:4]
  , input logic y
  , input tri1 logic jsiii [1:2][3:1]
  );
  
  
  nand ddfh(rry, oxexivok, iurbtodez);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   trireg logic [3:3][3:0]  iurbtodez -> logic iurbtodez
  
  not ipfuz(tqwijayyrr, oxexivok);
  
  not dvriyujbmz(ucdvac, y);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign tqwijayyrr = oxexivok;
  assign in = '{'{'b01,'b00x1}};
  assign iurbtodez = '{'{'b1,'b1zxz1,'b101z,'bz}};
  assign rry = 'b1;
  assign oxexivok = 'bz1;
endmodule: oqexmpwta

module ffedhkx
  ( output shortint ennhqb
  , output wire logic [0:2][1:4] lg [0:0][3:1][0:1][2:2]
  , output tri1 logic [3:3] k [4:2][3:0]
  , output realtime jed [2:4][4:0]
  , input shortreal eenai
  , input logic [3:0][4:1] uozyx [0:0][4:0]
  );
  
  wire logic [3:2] pczkrnxih [4:4];
  bit hk [2:1];
  tri1 logic wz [1:2][3:1];
  
  ptwxgn ivixh(.r(ngn), .qpzmph(hk), .bvuzha(atc), .twflb(eenai), .per(ennhqb), .mk(xqifqxg), .fpkakib(ennhqb));
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   trior logic [2:4]  r -> wire logic ngn
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:3][0:1][0:1][4:4]  bvuzha -> wire logic atc
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal eenai -> reg twflb
  //
  // warning: implicit conversion of port connection expands from 16 to 64 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint ennhqb -> time per
  //
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   wire logic xqifqxg -> logic [3:4][1:3]  mk
  //
  // warning: implicit conversion of port connection truncates from 16 to 9 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint ennhqb -> trior logic [0:2][2:4]  fpkakib
  
  xor tzyamjyc(ennhqb, ennhqb, ennhqb);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic ennhqb -> shortint ennhqb
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint ennhqb -> logic ennhqb
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   shortint ennhqb -> logic ennhqb
  
  oqexmpwta pys(.oxexivok(jr), .iurbtodez(vdyxojiyjq), .in(pczkrnxih), .y(eenai), .jsiii(wz));
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   trireg logic [3:3][3:0]  iurbtodez -> wire logic vdyxojiyjq
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal eenai -> logic y
  
  
  // Single-driven assigns
  assign jed = jed;
  
  // Multi-driven assigns
  assign atc = 'b10xzz;
  assign xqifqxg = ennhqb;
  assign wz = '{'{'b100x,'bx01x,'bz0x1},'{'b0101,'bx,'bxxxzz}};
  assign k = '{'{'{'b0z1x},'{'b000z},'{'bz00x0},'{'b0x}},'{'{'bzzx},'{'bzx1z0},'{'b0xzzz},'{'b1}},'{'{'bxzz},'{'bx},'{'b1xxz1},'{'b11x1x}}};
  assign lg = lg;
endmodule: ffedhkx



// Seed after: 15959535454375804453,5224943229413370507
