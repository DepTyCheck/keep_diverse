// Seed: 10640103557006565659,5224943229413370507

module u
  (input logic tfsnt [0:2][3:0], input tri0 logic cgoze [2:4][4:4], input logic [3:3][3:4][2:0]  utolhwivt);
  
  
  nand gstfmqkle(m, utolhwivt, utolhwivt);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [3:3][3:4][2:0]  utolhwivt -> logic utolhwivt
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  //   logic [3:3][3:4][2:0]  utolhwivt -> logic utolhwivt
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign cgoze = cgoze;
  assign m = 'bx0x0x;
endmodule: u

module hw
  ( output reg [0:0][0:4][3:0]  quzooinfe
  , output reg [4:2]  xnvl
  , output tri logic haa [0:3][1:3][3:3]
  , output supply1 logic [4:3] wbzasc [4:1][1:1][2:1]
  );
  
  
  not pcp(quzooinfe, quzooinfe);
  // warning: implicit conversion of port connection expands from 1 to 20 bits
  //   logic quzooinfe -> reg [0:0][0:4][3:0]  quzooinfe
  //
  // warning: implicit conversion of port connection truncates from 20 to 1 bits
  //   reg [0:0][0:4][3:0]  quzooinfe -> logic quzooinfe
  
  and wq(fevgt, xwrl, fevgt);
  
  
  // Single-driven assigns
  assign xnvl = '{'bz01,'bx0x00,'bzxx};
  
  // Multi-driven assigns
  assign haa = '{'{'{'bx0000},'{'b1},'{'b111}},'{'{'b1zx},'{'bz},'{'bxxz}},'{'{'b1},'{'bx},'{'b001z}},'{'{'b0zx00},'{'bzxzzz},'{'bzz}}};
endmodule: hw

module wqneddtxdr
  (input trior logic [0:0][2:2][0:1][2:0]  uo);
  
  tri0 logic mwbnk [2:4][4:4];
  logic zavlanvub [0:2][3:0];
  
  not kmu(ibs, wogudd);
  
  xor zpjasggsx(eevmaecf, eevmaecf, eevmaecf);
  
  u xi(.tfsnt(zavlanvub), .cgoze(mwbnk), .utolhwivt(wogudd));
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  //   wire logic wogudd -> logic [3:3][3:4][2:0]  utolhwivt
  
  
  // Single-driven assigns
  assign zavlanvub = zavlanvub;
  
  // Multi-driven assigns
  assign eevmaecf = 'bx01xz;
  assign mwbnk = mwbnk;
  assign wogudd = 'bx1z10;
endmodule: wqneddtxdr

module xadffomb
  (input logic [0:1][4:4][3:2] zdgf [1:0]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: xadffomb



// Seed after: 5678767469446421542,5224943229413370507
