// Seed: 3785318144795445061,5224943229413370507

module pqravuxwmh
  ( output wire logic acsow [1:1][2:1][1:3][4:4]
  , output wire logic [3:4][4:3][0:0][0:2] cjwc [0:2][3:0][1:2]
  , output logic sbyjznbx
  , output reg [2:1] xcnivan [1:3]
  );
  
  
  not vtii(bgpunmd, bgpunmd);
  
  and jrnuxjz(sbyjznbx, bgpunmd, y);
  
  nand l(xj, lnqw, kgqfljo);
  
  not emrym(bgpunmd, sbyjznbx);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kgqfljo = 'b1;
endmodule: pqravuxwmh

module v
  ( output longint g [1:0][1:3]
  , output supply0 logic [0:3][3:0][1:4][1:4]  s
  , input bit [2:4][1:2][0:4][2:0]  lhtoqzzst
  , input bit vpegann
  , input wire logic [3:1][2:4] tbsk [1:1][2:2]
  );
  
  
  nand ibrvwj(fb, s, lhtoqzzst);
  // warning: implicit conversion of port connection truncates from 256 to 1 bits
  //   supply0 logic [0:3][3:0][1:4][1:4]  s -> logic s
  //
  // warning: implicit conversion of port connection truncates from 90 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4][1:2][0:4][2:0]  lhtoqzzst -> logic lhtoqzzst
  
  
  // Single-driven assigns
  assign g = '{'{'b10,'b011,'b11110},'{'b0101,'b1,'b0}};
  
  // Multi-driven assigns
  assign s = '{'{'{'{'bx,'bzxz1,'b0z,'bx0x},'{'b00z0z,'bz,'bx00x,'b011zx},'{'bxzx,'b100,'bx,'b0},'{'b0,'b1,'b1z1,'b1xx}},'{'{'bx,'b11xx,'b11z,'b0zx1x},'{'bzx10,'bx,'b0x1,'b1},'{'bx,'b0,'b1,'b1xx1x},'{'b0z,'bxz,'b1x00x,'bzx}},'{'{'b0,'bzx,'b1x1,'b1z0},'{'bz0z0,'bz,'bx1z1,'b01},'{'b0zz,'b11,'bz00xx,'bxzxx},'{'b0z10,'b01x0x,'b11,'b001z}},'{'{'bzz1x,'b00x0x,'bxzx,'bzx1z1},'{'bxx1x,'bzz1x,'b11x,'b01xzz},'{'bz1z,'b1x,'b0,'b0xx},'{'b0,'b000,'b0z,'b10z11}}},'{'{'{'b0z0,'b0x01z,'b0z,'bzz},'{'b0100,'bxz00z,'bxxx,'bx1xx0},'{'bx,'b1,'bz,'b0xzx0},'{'bx,'b10,'bz1,'b0}},'{'{'b01011,'bz,'bx,'b11xz},'{'b10101,'bzxz,'b1,'b01},'{'b0x11,'bz1,'bx01,'b0z},'{'bx10z,'b1x,'b011,'bxz0}},'{'{'bx0xx,'b0z,'b1,'b11z},'{'bzz1xx,'bzz,'bx,'bxz},'{'bxzx,'b00,'b010z,'bz},'{'bz,'bxzx0z,'b101,'b10}},'{'{'bzz0z,'bz,'b01,'b0},'{'bz0,'bzz00,'bx1x0z,'b1},'{'b1,'bxz001,'bx1z0,'bz0},'{'b00110,'b1,'bz,'b100z1}}},'{'{'{'b0101x,'b0x1z,'bzz0zx,'bz011},'{'bx,'b0x1x,'bxz1,'bxx0},'{'bzzz0,'bzzzx,'bx,'b1},'{'b0x01,'b1z110,'bz0,'bzz1}},'{'{'bzz0zz,'bx0xzz,'bzxz1,'bx},'{'b0,'b01,'b0,'bx},'{'bzxx,'b11zxx,'bx0,'b00},'{'b11z0x,'b1x,'bxx,'b1x}},'{'{'b0,'bz,'bz,'b01},'{'b11xx,'b111,'bxxx,'bzzx},'{'b00z,'bz,'bx1z,'bz1z0},'{'bx110,'bz0,'b01zx,'b0z}},'{'{'bx0,'b11z,'b11xx0,'bx1},'{'bz00,'bxz,'bz0,'bxzz},'{'b1,'bzz0z,'bxx00x,'bxx},'{'bz1,'bz10,'b01,'b101xz}}},'{'{'{'bxx0,'bzzxx,'bz10,'b01},'{'b0z1x0,'bx,'b0xzx1,'bxzx1},'{'b0zxx,'bxxxx1,'bxxz,'bz01z},'{'bx,'b0x,'b110z,'bx0}},'{'{'bx,'bz1,'b01,'b01z01},'{'bx1zz,'bz0xx,'b11zzx,'b1z},'{'bzxx,'b0z,'bz1z,'bz00z1},'{'bx0zz1,'bzx00,'b0x1z,'b1}},'{'{'b1x,'bx1z10,'b1z101,'b00z},'{'bzx,'bzxx,'b0z,'bxx0},'{'b0,'b100zx,'bzzx1,'b01zzz},'{'bx1,'b1,'b0z1xz,'b0}},'{'{'b1z,'b1zxx,'b0x0,'b0},'{'b11,'bz,'b1z0,'bz01},'{'bzzz0,'b0,'bx,'b1z},'{'bxz,'bz,'b0x0,'bzx1xz}}}};
  assign tbsk = '{'{'{'{'bzx01,'bx1,'bxz},'{'b1x00,'bx0,'b0100},'{'bxxz0,'b1z100,'bz}}}};
  assign fb = 'b0xxz0;
endmodule: v

module uwgz
  ( output uwire logic [1:4][0:3] wbqilmwwz [3:1][1:4][4:3][4:4]
  , output bit [4:4][0:2]  tdhalkh
  , output trior logic [3:1][0:0] eixfpcci [2:2][1:2][0:1]
  , input logic [3:0]  vfabgutvyb
  , input logic unauap [1:0]
  , input longint rfjs [1:0]
  , input integer ereudagqkx [0:0]
  );
  
  
  nand ollmtfishj(smjd, tdhalkh, tdhalkh);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:2]  tdhalkh -> logic tdhalkh
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:2]  tdhalkh -> logic tdhalkh
  
  or hrzsoafcvk(a, tdhalkh, zs);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:2]  tdhalkh -> logic tdhalkh
  
  xor zdgc(ldhxsovbmg, tdhalkh, tdhalkh);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:2]  tdhalkh -> logic tdhalkh
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:4][0:2]  tdhalkh -> logic tdhalkh
  
  or yae(uxofarrh, ktmj, mosgrv);
  
  
  // Single-driven assigns
  assign wbqilmwwz = wbqilmwwz;
  assign tdhalkh = '{'{'b1010,'b101,'b0}};
  
  // Multi-driven assigns
  assign ldhxsovbmg = ldhxsovbmg;
  assign mosgrv = uxofarrh;
  assign ktmj = uxofarrh;
  assign eixfpcci = eixfpcci;
  assign zs = 'b01;
endmodule: uwgz



// Seed after: 911149662323965787,5224943229413370507
