// Seed: 4110387113029240658,5224943229413370507

module blliupw
  (output wire logic [3:0] utlywsc [2:2][0:4][3:3][4:2], output realtime ykxhynqx, input trireg logic [1:1]  gqodpwz);
  
  
  not zttwy(drjbbjctl, vzkfceh);
  
  not wj(gqodpwz, dltvlmnd);
  
  not djdr(b, wmwufd);
  
  or jv(egd, jbgxg, vzkfceh);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: blliupw

module uqp
  (output byte unnsjep);
  
  
  and z(rujd, ctldrl, rujd);
  
  nand pdunmrbq(unnsjep, unnsjep, ctldrl);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic unnsjep -> byte unnsjep
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte unnsjep -> logic unnsjep
  
  and h(ctldrl, grkugmggqv, unnsjep);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte unnsjep -> logic unnsjep
  
  not iopesqqtsv(eksb, grkugmggqv);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rujd = 'b011z0;
  assign eksb = 'b0x1;
  assign grkugmggqv = eksb;
  assign ctldrl = unnsjep;
endmodule: uqp



// Seed after: 13147908407365310562,5224943229413370507
