// Seed: 2626356992014929702,5224943229413370507

module llfxp
  ( output bit [0:2] umwkebxpy [0:2][3:3][0:0]
  , output wor logic [1:2][1:2][2:2] pfd [0:4][0:3][0:4]
  , input wand logic [3:2][0:0][2:1]  tq
  , input logic [0:2][4:4] vbvlsap [2:4]
  , input trireg logic [2:3][4:4][3:1][0:4] fgicbel [1:4][2:3]
  , input supply1 logic cphmpe [2:1][4:1]
  );
  
  
  not xowjv(bfhgtqfb, tq);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wand logic [3:2][0:0][2:1]  tq -> logic tq
  
  or uytmwnx(itusvbck, jngqunap, itusvbck);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign bfhgtqfb = 'bx100x;
  assign pfd = pfd;
endmodule: llfxp

module xzmin
  (output reg [2:0]  ilkzid);
  
  
  
  // Single-driven assigns
  assign ilkzid = ilkzid;
  
  // Multi-driven assigns
endmodule: xzmin

module igia
  ( output supply1 logic a [1:0]
  , output supply1 logic kcssmiy [1:0][1:1]
  , input bit [2:2][4:4] ni [2:3]
  , input logic [1:4][4:2]  ulhqvx
  , input reg xkvmaxj [0:4]
  , input tri1 logic [0:0][2:1][0:1]  tklhuaqrb
  );
  
  wor logic [1:2][1:2][2:2] utkejpqgzo [0:4][0:3][0:4];
  bit [0:2] wolryitcdf [0:2][3:3][0:0];
  supply1 logic arbcfxsyuo [2:1][4:1];
  trireg logic [2:3][4:4][3:1][0:4] lo [1:4][2:3];
  logic [0:2][4:4] vqtnrqbh [2:4];
  
  llfxp ardkhiz(.umwkebxpy(wolryitcdf), .pfd(utkejpqgzo), .tq(tklhuaqrb), .vbvlsap(vqtnrqbh), .fgicbel(lo), .cphmpe(arbcfxsyuo));
  
  and ogqyqvtb(wxdno, wxdno, lubws);
  
  not fvyfii(tklhuaqrb, txwx);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic tklhuaqrb -> tri1 logic [0:0][2:1][0:1]  tklhuaqrb
  
  nand tyiravk(tklhuaqrb, adwrdeemz, adwrdeemz);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic tklhuaqrb -> tri1 logic [0:0][2:1][0:1]  tklhuaqrb
  
  
  // Single-driven assigns
  assign vqtnrqbh = vqtnrqbh;
  
  // Multi-driven assigns
  assign arbcfxsyuo = arbcfxsyuo;
endmodule: igia



// Seed after: 7718581316640303111,5224943229413370507
