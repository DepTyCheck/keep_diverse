// Seed: 18330800851769687519,5224943229413370507

module ss
  (output realtime mnnqpxab, input tri0 logic [2:4][1:2][4:1] fnmw [1:4][1:0]);
  
  
  and vxrqsonijd(mgiobddvw, mnnqpxab, mnnqpxab);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime mnnqpxab -> logic mnnqpxab
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime mnnqpxab -> logic mnnqpxab
  
  not ai(mnnqpxab, mnnqpxab);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic mnnqpxab -> realtime mnnqpxab
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime mnnqpxab -> logic mnnqpxab
  
  and wem(zrfojn, e, e);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ss

module cpb
  ( output bit [1:0][1:2][3:4]  igapfoj
  , output wor logic [1:0] ynxyka [2:3][1:2][0:4][4:2]
  , output trior logic [0:1][1:0] qdckxsddk [0:3][1:0][0:3][1:4]
  , input reg [0:2][4:0][2:4]  iv
  , input wire logic [2:2][4:2] dp [3:1][4:3][0:1][4:0]
  , input time yq [0:2]
  , input trireg logic [2:3] hmalj [2:3][4:1][0:1]
  );
  
  
  
  // Single-driven assigns
  assign igapfoj = '{'{'{'b10,'b11100},'{'b01001,'b00}},'{'{'b11110,'b0011},'{'b0001,'b0}}};
  
  // Multi-driven assigns
  assign dp = dp;
  assign hmalj = '{'{'{'{'bz,'bxzxx},'{'bz1x,'bxx010}},'{'{'b1,'bz11},'{'b1z1xx,'bx1z}},'{'{'bxz,'b1x},'{'b00x,'b11z1x}},'{'{'bzxz0,'bz1},'{'bzz,'bz1}}},'{'{'{'bz1,'bxx11},'{'bzx0,'bxz}},'{'{'bxz110,'bxz},'{'b0x000,'b0x}},'{'{'bz10,'bz11},'{'b1xxx,'b0xz1}},'{'{'bx0,'bx0},'{'bx0,'b0xxx1}}}};
  assign ynxyka = ynxyka;
endmodule: cpb



// Seed after: 11249369895174539472,5224943229413370507
