// Seed: 31107661655320341,5224943229413370507

module i
  ( output reg oxlewkke
  , output logic [4:2][3:1][4:4][1:3]  mgj
  , input tri logic [1:1][1:1][4:2] lqywimfag [2:3]
  , input reg [1:3][2:1][0:1]  nwg
  );
  
  
  not vsjqed(bvuuiut, dgydnpiu);
  
  or vq(oa, oxlewkke, nwg);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [1:3][2:1][0:1]  nwg -> logic nwg
  
  
  // Single-driven assigns
  assign oxlewkke = 'bx00;
  
  // Multi-driven assigns
  assign dgydnpiu = oxlewkke;
  assign oa = 'bz0;
  assign bvuuiut = oxlewkke;
  assign lqywimfag = '{'{'{'{'b0z10z,'bx,'b0z1xz}}},'{'{'{'b1z0z1,'bz001,'b10}}}};
endmodule: i



// Seed after: 4328217436837865606,5224943229413370507
