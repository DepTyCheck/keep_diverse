// Seed: 5433596400001017772,5224943229413370507

module uzrjonz
  (output tri0 logic bxsbwqbpm [3:1][1:4][0:1][3:3], output wor logic [3:4][2:0][2:1][4:4] hkq [1:2], output logic [0:4][0:0]  v);
  
  
  not zrme(v, jhrqcpqjy);
  // warning: implicit conversion of port connection expands from 1 to 5 bits
  //   logic v -> logic [0:4][0:0]  v
  
  not bkdhtbrg(yuude, sseirzmcb);
  
  and znrogi(sseirzmcb, enyxqf, lccoch);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign lccoch = v;
endmodule: uzrjonz

module um
  (input reg [0:3][3:1][1:1]  fnleede);
  
  
  nand ob(jouhada, fnleede, jouhada);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [0:3][3:1][1:1]  fnleede -> logic fnleede
  
  not ke(yit, m);
  
  xor zrokocgmg(arkjgwnmce, m, fhj);
  
  not jtq(jouhada, fnleede);
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   reg [0:3][3:1][1:1]  fnleede -> logic fnleede
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign jouhada = yit;
  assign arkjgwnmce = 'bxzz;
  assign fhj = 'bz0z;
  assign m = 'bz01z;
  assign yit = 'bz0;
endmodule: um

module pmuzt
  ( output tri0 logic [3:2][1:2] rykw [2:4][0:0][2:0][4:3]
  , output reg [3:0][3:4]  hpplrm
  , output supply0 logic [0:3][2:4][3:3][4:2] mau [1:1][2:4]
  , output logic [2:0][3:3][4:1] ksyfijxt [4:1]
  , input trireg logic [1:0][0:2][0:2][1:2] uthhf [0:0][3:3]
  , input time rjiigyibj
  , input trireg logic [0:4]  pq
  , input supply0 logic v [0:0][4:0][2:4][0:1]
  );
  
  
  um lycbmm(.fnleede(rjiigyibj));
  // warning: implicit conversion of port connection truncates from 64 to 12 bits
  //   time rjiigyibj -> reg [0:3][3:1][1:1]  fnleede
  
  xor nxc(dugqypdb, hpplrm, pq);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  //   reg [3:0][3:4]  hpplrm -> logic hpplrm
  //
  // warning: implicit conversion of port connection truncates from 5 to 1 bits
  //   trireg logic [0:4]  pq -> logic pq
  
  um szjk(.fnleede(hpplrm));
  // warning: implicit conversion of port connection expands from 8 to 12 bits
  //   reg [3:0][3:4]  hpplrm -> reg [0:3][3:1][1:1]  fnleede
  
  not nokrqvnuk(hpplrm, cublimzcu);
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  //   logic hpplrm -> reg [3:0][3:4]  hpplrm
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: pmuzt

module bleg
  ( input wire logic [4:0][2:2][3:2][3:4] zlthq [3:0][3:3][1:0][1:3]
  , input bit [2:3][2:4][3:4][1:1]  euwn
  , input shortreal aockk
  , input realtime p
  );
  
  
  xor dwljzsyk(dpozcd, p, dpozcd);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime p -> logic p
  
  not s(dpozcd, p);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime p -> logic p
  
  not dlpsfhizf(ionblmesb, v);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign dpozcd = 'b1101;
  assign ionblmesb = dpozcd;
  assign v = 'b11zzx;
endmodule: bleg



// Seed after: 9771841626331172684,5224943229413370507
