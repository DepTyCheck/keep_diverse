// Seed: 3136145052316200612,5224943229413370507

module aalor
  (output reg [0:0][0:1][4:4] exomapjpw [2:4], input logic raosjk);
  
  
  nand rqj(ynvxhbo, zvy, ilcdmzrzgo);
  
  not tdluhu(x, ilcdmzrzgo);
  
  or kvajiaxt(zvy, ilcdmzrzgo, cijpul);
  
  
  // Single-driven assigns
  assign exomapjpw = '{'{'{'{'bx010x},'{'b10zz}}},'{'{'{'b0z},'{'bzx1x}}},'{'{'{'b11z0z},'{'bxx}}}};
  
  // Multi-driven assigns
  assign ynvxhbo = 'bz00;
  assign cijpul = zvy;
  assign zvy = ynvxhbo;
  assign ilcdmzrzgo = ynvxhbo;
endmodule: aalor



// Seed after: 8660179658830774611,5224943229413370507
