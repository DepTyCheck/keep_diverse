// Seed: 16902780496494233211,5224943229413370507

module rbz
  (input shortreal lgijbveav, input int nsoxmncw, input byte thmfiklf, input logic ydw);
  
  
  not hcnjg(dmogn, thmfiklf);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte thmfiklf -> logic thmfiklf
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: rbz

module mhaqylochf
  (input shortreal va [0:1][0:3], input supply0 logic uzr [0:1][1:1][0:1][3:1]);
  
  
  not bdqj(xpxdkkkb, ehsvnbp);
  
  or uvkfqfv(sqk, ehsvnbp, ehsvnbp);
  
  rbz l(.lgijbveav(ehsvnbp), .nsoxmncw(ehsvnbp), .thmfiklf(pikx), .ydw(ehsvnbp));
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic ehsvnbp -> shortreal lgijbveav
  //
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic ehsvnbp -> int nsoxmncw
  //
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic pikx -> byte thmfiklf
  
  or xhhstf(cpsegp, ehsvnbp, pikx);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xpxdkkkb = 'b1;
endmodule: mhaqylochf

module aitjf
  (output uwire logic [2:3] xhavblnr [0:1][1:4][3:4]);
  
  
  not n(lf, cxwifpro);
  
  nand cycd(cxwifpro, cxwifpro, cxwifpro);
  
  
  // Single-driven assigns
  assign xhavblnr = xhavblnr;
  
  // Multi-driven assigns
  assign cxwifpro = cxwifpro;
endmodule: aitjf

module oqizjm
  ( output wor logic [0:4][0:1][3:3][2:1] zd [1:3]
  , output real sfxeyxjbpj [3:4][0:2]
  , output logic [3:0][4:4]  ups
  , output supply1 logic [3:4] fypk [3:4]
  , input uwire logic [4:2][1:0] a [3:4][2:1][1:1]
  , input wand logic [2:4][2:3][3:1] ijnpeugo [0:0]
  , input reg [0:1][4:4] xowxwvdinl [3:2]
  , input reg [2:4] mrkithpw [0:2]
  );
  
  
  and am(pvpwcsmnx, ypeqolqa, ups);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   logic [3:0][4:4]  ups -> logic ups
  
  rbz cp(.lgijbveav(mcxlvcwqn), .nsoxmncw(alpb), .thmfiklf(ypeqolqa), .ydw(ups));
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic mcxlvcwqn -> shortreal lgijbveav
  //
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic alpb -> int nsoxmncw
  //
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wire logic ypeqolqa -> byte thmfiklf
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   logic [3:0][4:4]  ups -> logic ydw
  
  nand zrgvf(hhrybdwhsn, ups, ozhumdbvj);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   logic [3:0][4:4]  ups -> logic ups
  
  not s(ups, nj);
  // warning: implicit conversion of port connection expands from 1 to 4 bits
  //   logic ups -> logic [3:0][4:4]  ups
  
  
  // Single-driven assigns
  assign sfxeyxjbpj = '{'{'bz,'b1xxx,'b01x11},'{'bx,'b1100,'bz11}};
  
  // Multi-driven assigns
  assign zd = zd;
  assign pvpwcsmnx = nj;
  assign nj = ups;
  assign ypeqolqa = nj;
  assign fypk = fypk;
endmodule: oqizjm



// Seed after: 5024838802353150176,5224943229413370507
