// Seed: 17851572114395631375,5224943229413370507

module roshas
  ( output tri0 logic [2:2]  phduozjxn
  , output logic [2:2][0:0]  vvj
  , output tri1 logic [1:3][0:1] stnfvbd [1:2][3:3][2:4][1:4]
  , input logic [1:2][4:1][3:2]  miloydoyh
  , input tri logic [1:3][2:4][4:2][1:4] omfosnr [3:3][1:2]
  );
  
  
  
  // Single-driven assigns
  assign vvj = miloydoyh;
  
  // Multi-driven assigns
  assign phduozjxn = phduozjxn;
  assign omfosnr = omfosnr;
endmodule: roshas

module oycism
  (output bit [3:4] dol [2:3], input trior logic [3:1][3:2][2:4][3:4] nhegrbpq [4:3][0:1], input shortint dnzch [4:3][0:4]);
  
  
  not zgkcughhq(rkuo, wyrfydbb);
  
  not lblosbjdy(wyrfydbb, xjd);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign rkuo = wyrfydbb;
  assign nhegrbpq = nhegrbpq;
endmodule: oycism



// Seed after: 16778707474574903195,5224943229413370507
