// Seed: 8660179658830774611,5224943229413370507

module mbk
  (output supply1 logic [4:2][1:1][1:0] nf [4:4][0:1][1:2], output bit [3:2][1:1] udzbae [4:4][2:4]);
  
  
  
  // Single-driven assigns
  assign udzbae = udzbae;
  
  // Multi-driven assigns
  assign nf = nf;
endmodule: mbk

module f
  (output trior logic [3:0][4:1][0:0][2:1]  slwwojpj);
  
  
  xor xrlaaq(slwwojpj, slwwojpj, slwwojpj);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  //   logic slwwojpj -> trior logic [3:0][4:1][0:0][2:1]  slwwojpj
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  //   trior logic [3:0][4:1][0:0][2:1]  slwwojpj -> logic slwwojpj
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  //   trior logic [3:0][4:1][0:0][2:1]  slwwojpj -> logic slwwojpj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: f

module imiassfncp
  ( output tri logic [0:0][1:3] kdaffzin [4:2][2:0]
  , output bit [1:3][3:1][2:0][3:3]  taxfqzzhmb
  , output logic [2:4][2:1][0:4][4:3]  be
  , output reg [4:4][2:2] pbumi [3:4]
  , input time oscz
  , input supply0 logic [1:4][3:2][1:0] bfmbjtkf [3:0][0:2]
  , input tri0 logic rgisbektnd [3:1][4:3]
  );
  
  bit [3:2][1:1] ujufaoz [4:4][2:4];
  supply1 logic [4:2][1:1][1:0] t [4:4][0:1][1:2];
  
  not ncmouj(taxfqzzhmb, taxfqzzhmb);
  // warning: implicit conversion of port connection expands from 1 to 27 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic taxfqzzhmb -> bit [1:3][3:1][2:0][3:3]  taxfqzzhmb
  //
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:3][3:1][2:0][3:3]  taxfqzzhmb -> logic taxfqzzhmb
  
  mbk s(.nf(t), .udzbae(ujufaoz));
  
  or mq(be, taxfqzzhmb, taxfqzzhmb);
  // warning: implicit conversion of port connection expands from 1 to 60 bits
  //   logic be -> logic [2:4][2:1][0:4][4:3]  be
  //
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:3][3:1][2:0][3:3]  taxfqzzhmb -> logic taxfqzzhmb
  //
  // warning: implicit conversion of port connection truncates from 27 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:3][3:1][2:0][3:3]  taxfqzzhmb -> logic taxfqzzhmb
  
  not hm(symwnzkdt, be);
  // warning: implicit conversion of port connection truncates from 60 to 1 bits
  //   logic [2:4][2:1][0:4][4:3]  be -> logic be
  
  
  // Single-driven assigns
  assign pbumi = pbumi;
  
  // Multi-driven assigns
  assign bfmbjtkf = bfmbjtkf;
endmodule: imiassfncp



// Seed after: 16249125249849326094,5224943229413370507
