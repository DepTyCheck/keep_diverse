// Seed: 7679405928395605830,5224943229413370507

module mi
  (output wire logic [0:4][4:2] hpytk [0:2], input logic p, input supply0 logic [3:2][1:2]  lgeulj, input logic [3:3][2:1]  qvblo);
  
  
  not bkqutgzx(rhkqi, ripmon);
  
  nand ux(ripmon, ripmon, ripmon);
  
  not zjveoqkt(izqdaif, lgeulj);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   supply0 logic [3:2][1:2]  lgeulj -> logic lgeulj
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hpytk = hpytk;
  assign lgeulj = '{'{'bzz10,'b0z00},'{'bxz0z,'bxz1}};
  assign ripmon = 'b1x0;
endmodule: mi

module lhovg
  ( output trior logic [2:2][4:4][1:2][4:2] vg [0:3][1:1][3:2]
  , output triand logic [1:0][3:0][3:2]  ofwlxmz
  , output wor logic [3:2][3:0][0:1]  fk
  , output bit [2:0][0:4][2:3][1:4]  goeoqah
  , input tri logic [4:3][4:3] ffcargrzbk [3:4][1:1][0:4][2:0]
  , input bit [3:2][1:3] ofc [3:3][1:1]
  , input tri1 logic [3:4][2:4] rpjmc [2:0][0:0][1:0]
  , input triand logic [3:3][1:0] dlx [1:1][2:4][3:3][3:2]
  );
  
  
  nand oeu(goeoqah, jmkkpagv, nve);
  // warning: implicit conversion of port connection expands from 1 to 120 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic goeoqah -> bit [2:0][0:4][2:3][1:4]  goeoqah
  
  or cgwpizdm(buknnl, fk, rlkmgl);
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   wor logic [3:2][3:0][0:1]  fk -> logic fk
  
  or hjtrsdatxr(pbxdviqavs, pbxdviqavs, pbxdviqavs);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign pbxdviqavs = 'bz111;
endmodule: lhovg

module mkeygptij
  (output triand logic [1:2][0:3] evx [1:0], output real qvtnjkkq [0:3], output uwire logic [0:4][4:3][4:4][3:0] rrge [3:3]);
  
  trior logic [2:2][4:4][1:2][4:2] vywvjpn [0:3][1:1][3:2];
  triand logic [3:3][1:0] thiiltknm [1:1][2:4][3:3][3:2];
  tri1 logic [3:4][2:4] yg [2:0][0:0][1:0];
  bit [3:2][1:3] g [3:3][1:1];
  tri logic [4:3][4:3] hqp [3:4][1:1][0:4][2:0];
  
  not wbww(rksmzmtpx, qsusbmfqas);
  
  lhovg gzbepi(.vg(vywvjpn), .ofwlxmz(qsusbmfqas), .fk(qsusbmfqas), .goeoqah(xjx), .ffcargrzbk(hqp), .ofc(g), .rpjmc(yg), .dlx(thiiltknm));
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   triand logic [1:0][3:0][3:2]  ofwlxmz -> wire logic qsusbmfqas
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   wor logic [3:2][3:0][0:1]  fk -> wire logic qsusbmfqas
  //
  // warning: implicit conversion of port connection truncates from 120 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:0][0:4][2:3][1:4]  goeoqah -> wire logic xjx
  
  
  // Single-driven assigns
  assign rrge = rrge;
  assign g = g;
  assign qvtnjkkq = '{'b1,'bx,'b00xx,'bx0};
  
  // Multi-driven assigns
  assign thiiltknm = thiiltknm;
  assign qsusbmfqas = qsusbmfqas;
  assign evx = '{'{'{'b01x,'b10,'bxx1,'b1zx0},'{'bz01xx,'b0z,'bzz01,'bxxx0x}},'{'{'bxzzx,'bzxx1x,'bz,'b0x1x0},'{'bxzzzx,'bx0z,'bzz0z,'b1zx}}};
  assign rksmzmtpx = qsusbmfqas;
endmodule: mkeygptij

module hacdavklin
  ( input reg zsruokyru
  , input logic [4:0][0:4][1:4] ij [1:0]
  , input tri logic [0:3]  sckvzyq
  , input supply0 logic [4:3][0:3][4:1][2:2] pbjyyrra [4:2]
  );
  
  trior logic [2:2][4:4][1:2][4:2] edp [0:3][1:1][3:2];
  triand logic [3:3][1:0] obewhc [1:1][2:4][3:3][3:2];
  tri1 logic [3:4][2:4] mdrllkgjhu [2:0][0:0][1:0];
  bit [3:2][1:3] nezniwvyq [3:3][1:1];
  tri logic [4:3][4:3] h [3:4][1:1][0:4][2:0];
  
  lhovg r( .vg(edp)
         , .ofwlxmz(sckvzyq)
         , .fk(sckvzyq)
         , .goeoqah(ls)
         , .ffcargrzbk(h)
         , .ofc(nezniwvyq)
         , .rpjmc(mdrllkgjhu)
         , .dlx(obewhc)
         );
  // warning: implicit conversion of port connection truncates from 16 to 4 bits
  //   triand logic [1:0][3:0][3:2]  ofwlxmz -> tri logic [0:3]  sckvzyq
  //
  // warning: implicit conversion of port connection truncates from 16 to 4 bits
  //   wor logic [3:2][3:0][0:1]  fk -> tri logic [0:3]  sckvzyq
  //
  // warning: implicit conversion of port connection truncates from 120 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:0][0:4][2:3][1:4]  goeoqah -> wire logic ls
  
  
  // Single-driven assigns
  assign nezniwvyq = nezniwvyq;
  
  // Multi-driven assigns
  assign ls = zsruokyru;
  assign obewhc = obewhc;
  assign mdrllkgjhu = mdrllkgjhu;
  assign h = h;
endmodule: hacdavklin



// Seed after: 2232717311855488789,5224943229413370507
