// Seed: 18015104069983429213,5224943229413370507

module zoilqozltj
  ( output logic [0:3] uvu [3:2]
  , input realtime ebpfhbluh [1:2]
  , input reg zpaax [1:4]
  , input supply1 logic [4:3]  wsnnzfjbyd
  , input shortint evca
  );
  
  
  nand bzskn(ljlt, cdw, jns);
  
  not cvgjvsnng(cdw, cdw);
  
  nand eslxtx(mpwwkyj, lwj, jzhowunzci);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign cdw = 'b1zzx;
  assign lwj = wsnnzfjbyd;
  assign wsnnzfjbyd = cdw;
endmodule: zoilqozltj

module nkur
  (output tri1 logic zfbvgh [4:2][4:0][2:0], output reg [1:3][1:0]  ktoms);
  
  
  
  // Single-driven assigns
  assign ktoms = '{'{'b11z0,'bx1zz},'{'bxx,'b0},'{'bzzz,'bx1z0}};
  
  // Multi-driven assigns
  assign zfbvgh = '{'{'{'bxxzz,'b1111,'bzz1},'{'bzxz,'b0z111,'bx001},'{'b0x0,'b0xx11,'b0001},'{'b1z0z,'bx00x,'b1z1},'{'b1z1,'b00,'bxxzz}},'{'{'bz0,'b1,'bx0},'{'b10z1,'b10x,'bzx01},'{'bzz,'b0z1,'bz},'{'b10zz,'b0,'bz0},'{'b0,'bx1,'b1x00}},'{'{'b1x,'bz1000,'bxzzx},'{'bx1,'bz,'bz},'{'bx00zz,'bz,'b1},'{'b0zx0z,'b0,'bxx},'{'bz0,'bx,'bzxx}}};
endmodule: nkur



// Seed after: 16723051014337592514,5224943229413370507
