// Seed: 17257244788408976843,5224943229413370507

module ya
  ( output wand logic [2:0][0:0] ntibhmsvka [1:0][1:0][4:3][3:3]
  , output supply1 logic [1:4][0:1][0:0][2:3] pumk [2:2][0:1]
  , input realtime wokxpyed [4:1][0:0]
  , input bit [2:3][4:4] kfplp [4:1]
  , input wor logic [0:1][2:2][1:2][1:4] itcrkcw [2:4][4:3][4:0][1:0]
  , input reg [0:3][2:4][0:1][0:2]  actcvuk
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ntibhmsvka = ntibhmsvka;
endmodule: ya

module uyoq
  ( input tri logic [2:0][0:1][0:2] avfnkee [0:1][0:3][1:4]
  , input wand logic [0:2]  bjbozu
  , input logic m [2:3][0:2]
  , input longint vkutcln [4:2]
  );
  
  supply1 logic [1:4][0:1][0:0][2:3] deyles [2:2][0:1];
  wand logic [2:0][0:0] rbb [1:0][1:0][4:3][3:3];
  wor logic [0:1][2:2][1:2][1:4] uepnwm [2:4][4:3][4:0][1:0];
  bit [2:3][4:4] nigiyb [4:1];
  realtime ozwllnekv [4:1][0:0];
  
  or o(lfrqdwjtpz, tqjxc, tqjxc);
  
  ya owouddrt(.ntibhmsvka(rbb), .pumk(deyles), .wokxpyed(ozwllnekv), .kfplp(nigiyb), .itcrkcw(uepnwm), .actcvuk(tqjxc));
  // warning: implicit conversion of port connection expands from 1 to 72 bits
  //   wire logic tqjxc -> reg [0:3][2:4][0:1][0:2]  actcvuk
  
  
  // Single-driven assigns
  assign nigiyb = '{'{'{'b0000},'{'b0}},'{'{'b1},'{'b00010}},'{'{'b010},'{'b010}},'{'{'b01100},'{'b00110}}};
  assign ozwllnekv = ozwllnekv;
  
  // Multi-driven assigns
  assign rbb = rbb;
endmodule: uyoq

module bslmnkb
  ( output supply0 logic [4:1] uhbdcji [0:1]
  , output logic [0:2][3:2][3:4] wxvlhrgmqb [4:1]
  , output wor logic [4:2][2:0][2:0][3:4] rb [4:2]
  , input tri logic vi [0:4][2:1][4:0][4:2]
  , input tri logic [1:1][2:0]  iw
  , input supply1 logic [3:4][1:0][0:2][0:0] qbsoskcm [0:2][1:2]
  , input shortreal dhwx
  );
  
  
  and ghy(iw, iw, iw);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic iw -> tri logic [1:1][2:0]  iw
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri logic [1:1][2:0]  iw -> logic iw
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri logic [1:1][2:0]  iw -> logic iw
  
  or swk(iw, evigeswir, iw);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic iw -> tri logic [1:1][2:0]  iw
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri logic [1:1][2:0]  iw -> logic iw
  
  xor fwperlyde(kth, evigeswir, iw);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   tri logic [1:1][2:0]  iw -> logic iw
  
  
  // Single-driven assigns
  assign wxvlhrgmqb = '{'{'{'{'bzx10,'b111x},'{'bxzz,'b1}},'{'{'b11x0,'b1},'{'b0,'bz1}},'{'{'bz0xzz,'b0zxz},'{'b00000,'bxzxx}}},'{'{'{'bzx,'bzz},'{'bxx1,'bxx}},'{'{'b11z,'b0xz},'{'b10z01,'b0z001}},'{'{'b00,'bzxzz},'{'b1,'bz11x}}},'{'{'{'bx,'b0},'{'b11z1,'bz1x}},'{'{'bz00z1,'bzzx1},'{'bxzx01,'bzx00x}},'{'{'b0xz,'bz},'{'bxxx1,'b0}}},'{'{'{'b1110x,'bxxzx},'{'b0,'b0z11x}},'{'{'b11zx0,'b1},'{'bx,'b0z1}},'{'{'bx,'bz0xz1},'{'bx0xz,'b1}}}};
  
  // Multi-driven assigns
  assign uhbdcji = '{'{'bx,'bzxx,'b1xz,'b0x00},'{'bz,'b0x,'b00,'bxzx}};
  assign iw = '{'{'bx011,'b1,'b1xx0z}};
endmodule: bslmnkb



// Seed after: 8098496051366688625,5224943229413370507
