// Seed: 10771971825523251134,5224943229413370507

module zbukgdpt
  (output trior logic bgosrpdvre [0:4][2:0], output reg [4:2][1:2][4:4][1:0]  ixfagtiltq);
  
  
  
  // Single-driven assigns
  assign ixfagtiltq = '{'{'{'{'bx1z1,'b0}},'{'{'bz1z,'b11}}},'{'{'{'b010xz,'b0x001}},'{'{'b11z1z,'bx001}}},'{'{'{'b10100,'bzx0}},'{'{'bz,'bx1}}}};
  
  // Multi-driven assigns
  assign bgosrpdvre = '{'{'bx1,'b11x11,'bzx},'{'b1100,'bxxz1,'b1xz1},'{'bx11x1,'b00,'bzx01},'{'bx,'b0111,'b0x0x},'{'b10,'bx,'b0}};
endmodule: zbukgdpt

module k
  ( output tri0 logic [4:0][0:0][0:4][0:3]  ygfkdvsvm
  , output reg [4:0][1:3][3:3]  lxg
  , input reg gkjdaust
  , input bit [3:0][3:1] pkja [4:4]
  , input shortint u [4:0]
  );
  
  
  not fzu(ygfkdvsvm, iqjygf);
  // warning: implicit conversion of port connection expands from 1 to 100 bits
  //   logic ygfkdvsvm -> tri0 logic [4:0][0:0][0:4][0:3]  ygfkdvsvm
  
  xor ozkrrgya(ygfkdvsvm, lxg, lxg);
  // warning: implicit conversion of port connection expands from 1 to 100 bits
  //   logic ygfkdvsvm -> tri0 logic [4:0][0:0][0:4][0:3]  ygfkdvsvm
  //
  // warning: implicit conversion of port connection truncates from 15 to 1 bits
  //   reg [4:0][1:3][3:3]  lxg -> logic lxg
  //
  // warning: implicit conversion of port connection truncates from 15 to 1 bits
  //   reg [4:0][1:3][3:3]  lxg -> logic lxg
  
  xor exqw(ygfkdvsvm, hon, dynut);
  // warning: implicit conversion of port connection expands from 1 to 100 bits
  //   logic ygfkdvsvm -> tri0 logic [4:0][0:0][0:4][0:3]  ygfkdvsvm
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign hon = 'bz01;
endmodule: k



// Seed after: 12814626189442541259,5224943229413370507
