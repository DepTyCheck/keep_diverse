// Seed: 911149662323965787,5224943229413370507

module rhwmcjro
  (output integer zznol [3:4], input reg [1:3][3:2][2:3]  ytchgs, input bit [3:4][0:1][4:3][1:1]  vtbhi, input integer o);
  
  
  or jsfyegcobw(rakkynt, vtbhi, o);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:4][0:1][4:3][1:1]  vtbhi -> logic vtbhi
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   integer o -> logic o
  
  or zemcsvwfxx(hx, vtbhi, rakkynt);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:4][0:1][4:3][1:1]  vtbhi -> logic vtbhi
  
  not fgqtzycqyk(hx, wloi);
  
  xor xvc(udesyqndl, udesyqndl, vtbhi);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [3:4][0:1][4:3][1:1]  vtbhi -> logic vtbhi
  
  
  // Single-driven assigns
  assign zznol = zznol;
  
  // Multi-driven assigns
  assign wloi = vtbhi;
  assign hx = hx;
  assign udesyqndl = vtbhi;
  assign rakkynt = 'bz1110;
endmodule: rhwmcjro

module c
  (input logic cmcaxpp, input logic [2:3] hbzfagzjuh [4:2][4:3], input wor logic irkvirf);
  
  integer nvvl [3:4];
  
  rhwmcjro trjff(.zznol(nvvl), .ytchgs(cmcaxpp), .vtbhi(irkvirf), .o(cmcaxpp));
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic cmcaxpp -> reg [1:3][3:2][2:3]  ytchgs
  //
  // warning: implicit conversion of port connection expands from 1 to 8 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wor logic irkvirf -> bit [3:4][0:1][4:3][1:1]  vtbhi
  //
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic cmcaxpp -> integer o
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign irkvirf = irkvirf;
endmodule: c

module xibj
  ( input supply0 logic ytieo [2:4][3:0][2:1]
  , input realtime tjp
  , input wand logic [4:1][4:3][1:1] jbwjxgc [2:0][4:4][3:3]
  , input supply0 logic [4:2][3:1][2:2] najgiqjzby [2:4][3:0]
  );
  
  
  and v(igol, aqmeol, aqmeol);
  
  xor owmuq(vqfqkhob, igol, nkdjrqd);
  
  or a(aqmeol, nkdjrqd, tjp);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime tjp -> logic tjp
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign igol = aqmeol;
  assign nkdjrqd = aqmeol;
  assign aqmeol = tjp;
  assign ytieo = '{'{'{'b0,'bz1xz0},'{'b0z,'bx11z1},'{'b11z,'bz1x},'{'bz1,'b0z}},'{'{'b1zx,'b1z111},'{'bz0,'bx},'{'b110,'bzx10},'{'b1z,'b0x1}},'{'{'b101,'b0},'{'b10x,'b1z1},'{'bx,'b0110},'{'b0xz,'bxz}}};
  assign vqfqkhob = nkdjrqd;
endmodule: xibj

module alnqg
  (output wor logic [2:2][4:1][3:4] xvszcip [3:1][1:1][2:1][0:2], input reg [1:1][3:0]  t, input logic [4:0][3:4][1:2][4:2]  xibftn);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: alnqg



// Seed after: 1122856194526673955,5224943229413370507
