// Seed: 11791960886729708055,5224943229413370507

module yzxjprxvy
  ( output logic [3:1]  skavvptc
  , output reg [0:3]  onf
  , input tri0 logic [2:1] lqamtn [4:0]
  , input tri1 logic [0:4] gqqrskpjai [2:3][2:2][2:3][4:4]
  );
  
  
  not ovezdh(qhi, oedlgatsp);
  
  
  // Single-driven assigns
  assign skavvptc = onf;
  assign onf = skavvptc;
  
  // Multi-driven assigns
endmodule: yzxjprxvy

module eyrczbt
  (output tri logic yoc, output triand logic [4:1][4:1] cnnefag [2:0][2:3], output time unlzbrtj);
  
  
  or ipoxn(kojin, yoc, jobw);
  
  not c(cw, yoc);
  
  
  // Single-driven assigns
  assign unlzbrtj = yoc;
  
  // Multi-driven assigns
  assign jobw = yoc;
  assign cw = yoc;
  assign kojin = jobw;
  assign yoc = jobw;
  assign cnnefag = '{'{'{'{'b1x1,'b0z0,'bz0z1,'bz11zz},'{'b10z,'bzx10,'b10,'b0},'{'bx,'b10,'bx0x,'b1zx},'{'b01,'b1zz1x,'b11x,'b1x1}},'{'{'bxx11,'bx1xz,'b1,'b1},'{'b0xz,'b0x,'bz1x,'bz0x0},'{'b0,'bz,'bx1z,'bx},'{'b0z1x,'b1,'b0xzx,'b0}}},'{'{'{'bx0,'bzz11x,'b11z,'bz0zx},'{'bz1x,'bzz0,'bxxx10,'bz},'{'bx,'b1,'b0zz,'bz0z0},'{'b1z1,'bzzzz,'b0z0x,'bx1x0z}},'{'{'b111x,'bx0zz0,'b00,'bxxz},'{'bxx,'b1x0,'bz,'b1x},'{'bzx10,'bzx1,'b0010,'bxz1xz},'{'bz,'b0zzz,'b0110,'b1}}},'{'{'{'bz0,'bxx10,'bx1z0z,'b1101},'{'b0x,'b0z,'bz0z,'bx},'{'bz11z,'b1xx1x,'bx1x00,'bz},'{'bz,'b1111,'bzzzx,'bx0zz}},'{'{'bz0,'bz0,'bx,'b10010},'{'b0x11z,'bx,'bzx1z,'bz},'{'bx,'bz0,'bx1,'b01},'{'bx100z,'b1x1xx,'b1,'b01}}}};
endmodule: eyrczbt



// Seed after: 16166511167027967125,5224943229413370507
