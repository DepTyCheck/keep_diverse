// Seed: 10034344404040501477,5224943229413370507

module cswv
  (output shortreal p [1:3][2:3], input trireg logic kibjzunc [1:1]);
  
  
  not hfklxpbc(wamf, wamf);
  
  
  // Single-driven assigns
  assign p = '{'{'b1z11z,'bzzz},'{'b00x,'bzx1zz},'{'b01,'b00xx0}};
  
  // Multi-driven assigns
  assign wamf = 'bx1z;
  assign kibjzunc = '{'b000};
endmodule: cswv

module lbq
  (input bit [0:4][1:1] zjl [3:3], input integer znsvvwahd, input bit imwd [2:3], input uwire logic wgjzsuiwaa);
  
  
  and jbcvbbao(hmxjh, wgjzsuiwaa, wgjzsuiwaa);
  
  not qq(uasobprnyw, znsvvwahd);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   integer znsvvwahd -> logic znsvvwahd
  
  and vdjjaqsvxq(r, r, znsvvwahd);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   integer znsvvwahd -> logic znsvvwahd
  
  or qwioabtzbh(hmnrehefg, wgjzsuiwaa, hmnrehefg);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: lbq

module kymi
  ( output tri logic [4:2][2:4][4:3]  qflduf
  , output trior logic wcchgqvwl [4:1]
  , output supply1 logic [2:1][2:3] lic [1:1][4:4][2:1]
  , output bit zdush [2:1]
  );
  
  shortreal cqdnbqi [1:3][2:3];
  trireg logic ohyed [1:1];
  
  cswv a(.p(cqdnbqi), .kibjzunc(ohyed));
  
  
  // Single-driven assigns
  assign zdush = zdush;
  
  // Multi-driven assigns
  assign ohyed = '{'bxxz};
  assign lic = lic;
  assign wcchgqvwl = wcchgqvwl;
  assign qflduf = '{'{'{'bzxzz,'b1xx0},'{'bz1,'b1zx0z},'{'b10zx,'b00z}},'{'{'b0,'b1x},'{'b0,'b0xz},'{'bx1,'bz0}},'{'{'bzx1,'bxz},'{'bz0z0,'b1x0},'{'b10x1z,'b1zz1}}};
endmodule: kymi

module wrajiaadh
  ( output real yzrdia [3:0]
  , output supply1 logic [3:3][1:2]  edymvf
  , output wor logic [4:2][2:3][4:2][2:1] jhymviw [0:2][0:1]
  , input tri0 logic [2:0] wgqoch [4:2][4:3][0:1]
  , input supply0 logic [0:1][1:0][0:0][1:1] ayoggx [2:1]
  , input shortint ivdq [4:0]
  );
  
  bit kpablmh [2:1];
  supply1 logic [2:1][2:3] aj [1:1][4:4][2:1];
  trior logic mctrx [4:1];
  
  or gzo(musiwtgx, edymvf, musiwtgx);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   supply1 logic [3:3][1:2]  edymvf -> logic edymvf
  
  kymi arudycmxij(.qflduf(edymvf), .wcchgqvwl(mctrx), .lic(aj), .zdush(kpablmh));
  // warning: implicit conversion of port connection truncates from 18 to 2 bits
  //   tri logic [4:2][2:4][4:3]  qflduf -> supply1 logic [3:3][1:2]  edymvf
  
  
  // Single-driven assigns
  assign yzrdia = yzrdia;
  
  // Multi-driven assigns
  assign edymvf = '{'{'b00x,'bx1z10}};
  assign wgqoch = '{'{'{'{'bz0,'b110,'b0},'{'b11z1,'b1z10z,'bxz1}},'{'{'b1,'bzx00,'bx1x},'{'bx10,'b010zz,'b1xxz}}},'{'{'{'bz,'bzz0,'b0},'{'b1z,'b0z11,'bx}},'{'{'bzz1,'bz,'b0z0},'{'bz10zx,'b11,'bx}}},'{'{'{'bxz1z1,'b110,'b00},'{'bz,'bxxz,'b11x0}},'{'{'b1x010,'b11,'b01},'{'bz0,'bx10,'b1}}}};
  assign ayoggx = ayoggx;
  assign musiwtgx = musiwtgx;
  assign jhymviw = jhymviw;
endmodule: wrajiaadh



// Seed after: 6347729663862269036,5224943229413370507
