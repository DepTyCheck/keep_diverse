// Seed: 12034918165399613485,5224943229413370507

module tiyzfk
  ( output triand logic [4:4][4:3][1:2] nm [2:3][2:1][0:0][2:1]
  , output realtime mhxfnn
  , output bit [0:2][1:2]  wqshkch
  , input integer dcx
  , input logic [4:4][1:2][1:0]  gaj
  , input uwire logic aabma
  );
  
  
  xor gupt(qm, mhxfnn, dcx);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime mhxfnn -> logic mhxfnn
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   integer dcx -> logic dcx
  
  and vad(hhjlbmqta, wqshkch, aabma);
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:2][1:2]  wqshkch -> logic wqshkch
  
  not wo(wqshkch, mhxfnn);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic wqshkch -> bit [0:2][1:2]  wqshkch
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime mhxfnn -> logic mhxfnn
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: tiyzfk

module nwhzfvul
  ( output bit [1:2][3:0][2:1]  zkewfa
  , output wire logic pwnghsqeo [0:0][4:3][3:1][1:2]
  , output bit [4:4][3:3]  pqsjolpf
  , output trior logic [3:3] pgulzk [0:3][1:4][3:4][4:0]
  );
  
  
  not qbwrz(zkewfa, jveg);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic zkewfa -> bit [1:2][3:0][2:1]  zkewfa
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign pwnghsqeo = '{'{'{'{'bx0z,'b011},'{'bxz0,'b01z0z},'{'bxxz,'b1}},'{'{'b001x,'bz},'{'bz,'bx1z0z},'{'b1z0,'bxzz}}}};
endmodule: nwhzfvul



// Seed after: 16188638392432509924,5224943229413370507
