// Seed: 15853465871684603681,5224943229413370507

module nndz
  ( output reg gikybab [3:4][1:3]
  , output tri logic [2:2][1:0][3:1][1:4] ads [4:3][2:2][1:4][2:0]
  , output reg [3:1][0:1]  ewgtcyo
  , output reg wozozd
  );
  
  
  xor mnyyl(ieomac, wozozd, a);
  
  not wfveeqxqb(w, kk);
  
  not nbkvwtizya(kk, xhi);
  
  
  // Single-driven assigns
  assign gikybab = '{'{'b1zx,'bx00,'b0011},'{'bxx110,'bz001x,'b1z1z}};
  assign wozozd = xhi;
  assign ewgtcyo = ewgtcyo;
  
  // Multi-driven assigns
  assign xhi = ieomac;
  assign a = 'bx1x;
  assign ads = ads;
  assign ieomac = kk;
  assign w = 'bx0zz0;
endmodule: nndz



// Seed after: 2097695163638439650,5224943229413370507
