// Seed: 12515504994790153200,5224943229413370507

module mmvvhyzzuh
  ( output bit stbtx [2:1][4:4]
  , output reg [2:4][1:1]  j
  , output bit [4:4][3:4]  gl
  , output trior logic [4:1] wdbzhk [2:3]
  , input tri logic paxuigj [1:1][2:3]
  , input int guace
  , input bit wqgcww
  , input tri logic [0:2][0:0][4:0]  yznydxfp
  );
  
  
  not hbuywcj(j, wqgcww);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic j -> reg [2:4][1:1]  j
  //
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit wqgcww -> logic wqgcww
  
  
  // Single-driven assigns
  assign stbtx = '{'{'b000},'{'b0}};
  assign gl = '{'{'b01,'b0}};
  
  // Multi-driven assigns
  assign wdbzhk = wdbzhk;
endmodule: mmvvhyzzuh

module gcsz
  ( output shortreal pjj [3:2][4:4]
  , output tri0 logic [3:0] pccmcvlulm [2:0][2:1][4:3]
  , input wire logic [3:3][0:0][3:0] unjevswql [1:2][1:1][2:3][3:2]
  );
  
  
  not pocuvj(dnzcyw, cdonyswte);
  
  not apjnyr(xbuaxmj, hxhym);
  
  
  // Single-driven assigns
  assign pjj = '{'{'b0110x},'{'bx}};
  
  // Multi-driven assigns
  assign unjevswql = unjevswql;
endmodule: gcsz

module hxczkzclb
  ( output wand logic [0:1][4:3] fwncomsmyj [3:4][2:0][3:3][4:3]
  , input reg [0:2]  eoerbbjdds
  , input supply0 logic fbq [3:1]
  , input tri0 logic [0:4][2:0] eieuaht [1:1][3:1]
  , input wire logic [4:4] nmxwordydl [2:1][4:2][0:3][3:0]
  );
  
  tri0 logic [3:0] jtgmb [2:0][2:1][4:3];
  shortreal oqcvdsnqiv [3:2][4:4];
  wire logic [3:3][0:0][3:0] rmjkfmytmq [1:2][1:1][2:3][3:2];
  
  and oclc(digcosnkgi, oozwnm, oozwnm);
  
  not qlstkjft(mvmscfmf, ahro);
  
  gcsz racy(.pjj(oqcvdsnqiv), .pccmcvlulm(jtgmb), .unjevswql(rmjkfmytmq));
  
  not vq(wshkaf, zyxikblhjb);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign eieuaht = '{'{'{'{'bzz001,'bxz0,'bx},'{'b1,'b00xx0,'bzz1},'{'bzx0,'bzz,'b0x},'{'bzzx,'b001,'b1},'{'bzz1z,'b1010,'b10x0}},'{'{'b00,'bxx,'b00},'{'b00xz1,'bz101,'bz1zzx},'{'b11,'b11xz1,'b0},'{'b1xzz,'b011,'b1},'{'b10,'b0xzx,'b0x0xx}},'{'{'bx,'bzx01,'b0x00},'{'bz010x,'bzx1x,'bzx1},'{'bx01,'b1x1,'b111x},'{'bx1xz,'bz,'b10z},'{'bzz0xx,'b00,'b1x}}}};
  assign jtgmb = '{'{'{'{'bx00,'b0x,'b11x,'b1x1z},'{'bxzx,'b1z1z,'b11x,'bx}},'{'{'b0z1xx,'bxxx1x,'bx,'b01},'{'b01z1,'bx,'b0z,'b1z11x}}},'{'{'{'bz1zz,'bxz10,'b00,'b1},'{'b0x,'b11,'b11x0x,'b0}},'{'{'b00xz,'b1z00,'b0011x,'bzzx1},'{'b1,'b1,'bz0x,'bzz}}},'{'{'{'b1z0x1,'bx,'b01,'b0},'{'bxz1,'bx1x,'b1,'b1z0zx}},'{'{'b111,'b01x0z,'bzx1,'b0zz0},'{'b1,'b0x,'b10z1x,'bz101}}}};
  assign oozwnm = zyxikblhjb;
  assign zyxikblhjb = 'bx001z;
  assign fwncomsmyj = fwncomsmyj;
endmodule: hxczkzclb



// Seed after: 17194071564510378098,5224943229413370507
