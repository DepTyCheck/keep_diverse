// Seed: 16058725124331033669,5224943229413370507

module uengql
  (output reg [2:0][4:2]  eqx, output wand logic [1:3][3:3]  eqy, output bit [1:4][3:3][0:2]  upykuqt, output real pu);
  
  
  not msdidqi(whgeridh, eqx);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  //   reg [2:0][4:2]  eqx -> logic eqx
  
  and cztaeka(pu, rxvvvr, eqy);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic pu -> real pu
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   wand logic [1:3][3:3]  eqy -> logic eqy
  
  
  // Single-driven assigns
  assign eqx = '{'{'b0z,'bxz0,'bz0},'{'bx1x,'b0,'bx0},'{'b10x,'b11,'bxx10}};
  assign upykuqt = '{'{'{'b10010,'b0111,'b1111}},'{'{'b1,'b0110,'b11}},'{'{'b01111,'b1011,'b10}},'{'{'b0,'b0,'b00}}};
  
  // Multi-driven assigns
  assign rxvvvr = 'b11z00;
  assign eqy = eqx;
  assign whgeridh = 'bz1z;
endmodule: uengql

module jvopmdcsh
  (output longint okgfddepg);
  
  
  uengql outz(.eqx(ehjnbk), .eqy(okgfddepg), .upykuqt(w), .pu(yiuxbjvh));
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  //   reg [2:0][4:2]  eqx -> wire logic ehjnbk
  //
  // warning: implicit conversion of port connection expands from 3 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   wand logic [1:3][3:3]  eqy -> longint okgfddepg
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [1:4][3:3][0:2]  upykuqt -> wire logic w
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   real pu -> wire logic yiuxbjvh
  
  not pbp(w, w);
  
  not imoehno(yiuxbjvh, ehjnbk);
  
  not uhxblm(yiuxbjvh, gv);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign w = okgfddepg;
  assign yiuxbjvh = ehjnbk;
  assign gv = okgfddepg;
  assign ehjnbk = w;
endmodule: jvopmdcsh



// Seed after: 1250704759608574705,5224943229413370507
