// Seed: 8101242052950840334,5224943229413370507

module cldozwif
  ( output logic [4:4][4:0][4:0][4:0]  mrseodlzhl
  , output reg fghs
  , output longint gawc
  , input wire logic vttxuem [3:0]
  , input logic lfpjl
  );
  
  
  
  // Single-driven assigns
  assign gawc = mrseodlzhl;
  assign fghs = mrseodlzhl;
  assign mrseodlzhl = mrseodlzhl;
  
  // Multi-driven assigns
  assign vttxuem = '{'bx10,'bx,'bzzx0,'b0x100};
endmodule: cldozwif

module jjubsk
  (output logic [4:1][3:4][1:1] ddquv [4:0], input wor logic [1:2] zibto [1:1][4:4][3:2][1:3]);
  
  
  not jwni(aogcvqc, an);
  
  not yft(dsmitze, an);
  
  nand ypbopenq(an, qvlbaj, iejzowvxc);
  
  not azjfi(hz, nnopkvjtg);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: jjubsk

module yqxt
  ( output logic [3:3][4:1][0:2] ky [2:3]
  , output shortreal oxbu [3:3][0:0]
  , output supply1 logic [3:2][2:4] hvbevfsuq [4:0][0:0][0:1][4:3]
  , input supply1 logic [0:2][3:0][4:4][2:3] xyhs [4:2][4:1][3:0]
  , input tri logic [1:2][1:1] cvipmteu [2:0][4:1][3:0][3:0]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign xyhs = xyhs;
  assign cvipmteu = cvipmteu;
endmodule: yqxt

module jrrjzpk
  (output reg [3:0][2:2][2:4][4:1]  xub);
  
  logic [4:1][3:4][1:1] plsyrhlk [4:0];
  wor logic [1:2] avezwe [1:1][4:4][3:2][1:3];
  
  not aja(oucoodsp, c);
  
  jjubsk lxukms(.ddquv(plsyrhlk), .zibto(avezwe));
  
  nand eshuet(hjstwh, c, c);
  
  not akjy(xub, c);
  // warning: implicit conversion of port connection expands from 1 to 48 bits
  //   logic xub -> reg [3:0][2:2][2:4][4:1]  xub
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: jrrjzpk



// Seed after: 15475924140465045634,5224943229413370507
