// Seed: 9916430053765975954,5224943229413370507

module tfxczjy
  (output trior logic [1:3] yoemqv [2:0][3:1][2:4][1:0], input trior logic njejkuo [0:1][3:0][1:4][4:3]);
  
  
  not kvzadaod(rsaljcdnfc, rsaljcdnfc);
  
  not yf(fu, oxoasikb);
  
  not rlamtmi(drnuteb, z);
  
  nand ogrnnrjedo(drnuteb, rsaljcdnfc, v);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign yoemqv = yoemqv;
  assign z = rsaljcdnfc;
  assign rsaljcdnfc = rsaljcdnfc;
  assign fu = fu;
  assign njejkuo = '{'{'{'{'bx,'bx},'{'b0,'b1},'{'b0z,'b11001},'{'bz,'bx0x}},'{'{'b1,'b01xzz},'{'b000,'b00z},'{'bxzxzz,'bx00},'{'bxz11x,'b1x0}},'{'{'b0,'bx1x},'{'b0,'bx11z},'{'b0z,'bx010},'{'bxzz0,'b0}},'{'{'b0z,'b11010},'{'bx0xzx,'b1xz1x},'{'bx,'bx1xz0},'{'b10,'b01zxz}}},'{'{'{'b100,'bz},'{'bzz,'b0010x},'{'bzz,'bx},'{'bx10,'b1}},'{'{'b0zzxx,'b110},'{'bz0xx,'b01},'{'bx,'b1z0},'{'bz0x,'b0101}},'{'{'b01,'bzz0},'{'bzx,'bx},'{'b111x,'bx},'{'b1x00,'b10}},'{'{'b100,'b0},'{'b1,'b0x1},'{'b1,'bx11},'{'bx0,'bzx0}}}};
endmodule: tfxczjy

module pzzuwps
  ( output logic [0:2][4:4]  cedgmfvh
  , output logic [2:1][3:1] iqatyyhvpj [1:0]
  , output tri1 logic amlnselp [3:2][4:2][4:4][4:3]
  , output tri1 logic [4:1][0:4][3:4] ulgxu [0:2]
  , input time kigow
  , input uwire logic [1:1][3:1][0:3] ffnfzmtif [3:3]
  , input wand logic vfmctk [4:2][0:3][2:0][0:2]
  , input trior logic [0:1][0:1][0:4] caxwrfay [4:2][1:2]
  );
  
  trior logic [1:3] imxop [2:0][3:1][2:4][1:0];
  trior logic [1:3] gyvqcp [2:0][3:1][2:4][1:0];
  trior logic jz [0:1][3:0][1:4][4:3];
  
  tfxczjy um(.yoemqv(gyvqcp), .njejkuo(jz));
  
  xor c(gewknid, gmpurdypt, cedgmfvh);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   logic [0:2][4:4]  cedgmfvh -> logic cedgmfvh
  
  tfxczjy mhyayvgftn(.yoemqv(imxop), .njejkuo(jz));
  
  xor qaptrez(cedgmfvh, gmpurdypt, cedgmfvh);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic cedgmfvh -> logic [0:2][4:4]  cedgmfvh
  //
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  //   logic [0:2][4:4]  cedgmfvh -> logic cedgmfvh
  
  
  // Single-driven assigns
  assign iqatyyhvpj = '{'{'{'b1zzzx,'bz11z,'bxxzz1},'{'bx101,'b10,'bxx11}},'{'{'bx,'b11z01,'bz1},'{'bx01,'bx11zz,'b0z10}}};
  
  // Multi-driven assigns
  assign gmpurdypt = 'b1zz;
  assign caxwrfay = caxwrfay;
  assign jz = '{'{'{'{'b0z,'b01z01},'{'bxz1,'b0},'{'b0z0x,'b0z},'{'bx0,'b010}},'{'{'b0zz,'bz},'{'b11x,'b0x},'{'b0,'b11z11},'{'bx01,'b0x0z}},'{'{'b10x,'b1},'{'b00,'b10},'{'b1000z,'b0x1},'{'b1,'b0z}},'{'{'b0zz01,'bz},'{'bzx1x,'bxz111},'{'bz0,'b00z01},'{'bzz0z,'b00z10}}},'{'{'{'b1xz1,'b10},'{'bzz11,'b01},'{'b0,'b11z},'{'bx000,'bxx0}},'{'{'b1z,'bx00z},'{'b111,'bx},'{'b1xzxx,'b1z1},'{'bzx,'bz}},'{'{'bz100,'bxzz0},'{'bz,'b0xx},'{'b01x,'b0z1},'{'b0,'bx1xz1}},'{'{'b00x0x,'bz0z},'{'bz0x1,'b11x0z},'{'b1x00z,'b100x},'{'b0zx,'b0z0z}}}};
  assign ulgxu = ulgxu;
  assign amlnselp = '{'{'{'{'bx,'bx}},'{'{'bzxx1,'bz0x01}},'{'{'bzz0,'b11x}}},'{'{'{'bx0x0,'bzz}},'{'{'bz,'b0x11}},'{'{'bxz0z1,'bzxz0}}}};
endmodule: pzzuwps



// Seed after: 8288159748330704549,5224943229413370507
