// Seed: 2097695163638439650,5224943229413370507

module zhbw
  ( input logic [2:3][2:4][4:2]  adhljqjidc
  , input shortint htpek
  , input tri0 logic liiau [3:0][2:2][4:0]
  , input wor logic [1:3] ubq [2:3][4:1][3:0][2:3]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign liiau = liiau;
  assign ubq = ubq;
endmodule: zhbw



// Seed after: 13898922656242679089,5224943229413370507
