// Seed: 8098496051366688625,5224943229413370507

module rqigpys
  ( output tri1 logic [4:2][0:3][0:0][1:3] x [3:2][4:4]
  , output uwire logic tx
  , output wor logic [0:0]  rzgju
  , output wor logic [4:3][1:1][3:1][1:1] yyhof [2:0]
  , input realtime hwiequky
  );
  
  
  xor aeeaynhnyn(aefarjtxx, rwco, tx);
  
  not cjijry(znpeb, rwco);
  
  nand xas(erwcqivwbe, rzgju, jcozxltrhe);
  
  not e(dw, tx);
  
  
  // Single-driven assigns
  assign tx = 'bzz;
  
  // Multi-driven assigns
  assign erwcqivwbe = 'bzz;
  assign znpeb = tx;
  assign x = x;
endmodule: rqigpys

module sirx
  (output reg bamtemjrcf [2:3], input wand logic [2:4][3:2][0:1][3:2]  gvkrzpb, input tri0 logic [1:1] lmnnjqwczz [2:0][0:4]);
  
  wor logic [4:3][1:1][3:1][1:1] p [2:0];
  tri1 logic [4:2][0:3][0:0][1:3] ss [3:2][4:4];
  
  rqigpys pacw(.x(ss), .tx(grua), .rzgju(gvkrzpb), .yyhof(p), .hwiequky(gvkrzpb));
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   wor logic [0:0]  rzgju -> wand logic [2:4][3:2][0:1][3:2]  gvkrzpb
  //
  // warning: implicit conversion of port connection expands from 24 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wand logic [2:4][3:2][0:1][3:2]  gvkrzpb -> realtime hwiequky
  
  not kwpsvt(ojdl, gvkrzpb);
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   wand logic [2:4][3:2][0:1][3:2]  gvkrzpb -> logic gvkrzpb
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign p = p;
  assign ss = ss;
  assign gvkrzpb = '{'{'{'{'bx111z,'bxz},'{'bzxzz0,'bz0xzx}},'{'{'bx10z,'b1},'{'b1z,'bxzx10}}},'{'{'{'bzx,'bzxz1x},'{'bz11xx,'bxxx10}},'{'{'bx0z1x,'b0z111},'{'bzzx0x,'b01z}}},'{'{'{'bzx,'b1xxzz},'{'bxxzz1,'bxz}},'{'{'bzz0,'bzz0},'{'bz,'b0z}}}};
  assign ojdl = gvkrzpb;
endmodule: sirx

module eobw
  ( output trireg logic [1:3] mzgdmnv [2:3][2:1][0:2]
  , output reg [3:1][4:4] v [1:1]
  , input uwire logic wnvq [1:3][2:1][2:2]
  , input reg [3:1][0:2]  jpja
  , input logic y [3:4]
  , input logic mnhcudtrrx
  );
  
  wor logic [4:3][1:1][3:1][1:1] rtmnpkz [2:0];
  tri1 logic [4:2][0:3][0:0][1:3] ipnzhlfsyu [3:2][4:4];
  reg axxuppq [2:3];
  tri0 logic [1:1] s [2:0][0:4];
  
  nand xdt(cizjsnctrz, mnhcudtrrx, mnhcudtrrx);
  
  or pe(beavzb, beavzb, mnhcudtrrx);
  
  sirx ejp(.bamtemjrcf(axxuppq), .gvkrzpb(mnhcudtrrx), .lmnnjqwczz(s));
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   logic mnhcudtrrx -> wand logic [2:4][3:2][0:1][3:2]  gvkrzpb
  
  rqigpys eemexevscp(.x(ipnzhlfsyu), .tx(beavzb), .rzgju(ycv), .yyhof(rtmnpkz), .hwiequky(beavzb));
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   wire logic beavzb -> realtime hwiequky
  
  
  // Single-driven assigns
  assign v = '{'{'{'bx},'{'b1},'{'b1zz0}}};
  
  // Multi-driven assigns
  assign ycv = 'b0x0;
endmodule: eobw

module ehnrjmtfu
  ( output logic [2:2]  baijdzfb
  , input shortreal vnumhhjr [4:0][4:4][0:1]
  , input supply0 logic [0:0][3:1][1:4] svqqlv [2:1][2:2]
  , input bit [0:2][1:3][1:0]  wybkgn
  );
  
  
  
  // Single-driven assigns
  assign baijdzfb = '{'b001};
  
  // Multi-driven assigns
  assign svqqlv = svqqlv;
endmodule: ehnrjmtfu



// Seed after: 1913518407355023998,5224943229413370507
