// Seed: 17194071564510378098,5224943229413370507

module th
  ( output reg [4:2]  norbhub
  , output reg [1:3][2:0][1:1] lr [0:1]
  , input tri0 logic [4:0] ifloksfak [4:2]
  , input bit kbekaxfn [0:0]
  , input reg [2:4] icple [2:1][2:0][2:0]
  , input wand logic [4:2][1:1] wgujxv [4:3][2:2][4:2][0:4]
  );
  
  
  
  // Single-driven assigns
  assign norbhub = norbhub;
  assign lr = lr;
  
  // Multi-driven assigns
  assign ifloksfak = ifloksfak;
  assign wgujxv = wgujxv;
endmodule: th



// Seed after: 7679405928395605830,5224943229413370507
