// Seed: 15959535454375804453,5224943229413370507

module gsk
  (output byte lstwc [3:0][4:2], input logic [2:0][4:4][3:0]  c);
  
  
  and odgamnd(uxwsxqcwiw, hzle, hxzs);
  
  nand xxlcjouzd(hzle, hxzs, ahrqfdtqzh);
  
  not r(hzle, gr);
  
  nand kjwkxgfi(iznjlpa, hzle, ahrqfdtqzh);
  
  
  // Single-driven assigns
  assign lstwc = lstwc;
  
  // Multi-driven assigns
  assign hzle = 'b1zx00;
  assign gr = c;
  assign ahrqfdtqzh = 'bzzz00;
  assign iznjlpa = 'b0;
  assign hxzs = 'b001x0;
endmodule: gsk

module sdtsbox
  ( output wire logic [1:2][0:4][1:4][1:2] v [0:3][2:1]
  , input bit [1:1][3:0][3:2][0:1]  grfmbinv
  , input supply0 logic [4:3][0:2][0:3][0:3] rpusywp [0:4][3:4][3:1][3:2]
  , input bit [3:3][2:1][2:3] fkhrh [2:3]
  );
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign v = v;
  assign rpusywp = rpusywp;
endmodule: sdtsbox

module vktbhtubeo
  (input reg [2:4] qakjoqni [4:0], input reg aoglrebres, input realtime c, input tri0 logic [4:2][4:2][2:2] kbaoim [0:0]);
  
  
  nand zky(rvwfepbh, ynoowsv, c);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime c -> logic c
  
  not gmewumjimy(ynoowsv, alp);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign alp = ynoowsv;
endmodule: vktbhtubeo

module i
  ( output triand logic [4:2][0:2][3:2] gax [4:4][1:4][2:4][1:4]
  , output triand logic [3:4][1:4] twvfgxiur [1:0][4:2][1:2][0:1]
  , output logic [2:4][0:3][0:4]  uvehixhwth
  , output wire logic [1:2][1:0][1:2] bciqvya [3:0]
  );
  
  
  
  // Single-driven assigns
  assign uvehixhwth = uvehixhwth;
  
  // Multi-driven assigns
  assign gax = gax;
  assign bciqvya = '{'{'{'{'b1x1,'bz1},'{'b11x,'b1x1}},'{'{'bx0,'b1z1},'{'b1x10z,'b11}}},'{'{'{'b00,'bx},'{'b10,'bz011}},'{'{'bz,'b0z101},'{'bx1z00,'b100x}}},'{'{'{'b111,'b00z},'{'b0xx,'bx11z}},'{'{'bx10z,'bzx1x},'{'b101,'bz11z0}}},'{'{'{'b0,'bzz1xx},'{'bx011z,'bxx0}},'{'{'bxxx0,'bz1},'{'b1z11,'b0101x}}}};
endmodule: i



// Seed after: 3807221459878586453,5224943229413370507
