// Seed: 7587504049292560125,5224943229413370507

module zb
  (output trireg logic [1:2][2:3] qtqmqrax [2:3][2:4][1:4][4:1]);
  
  
  nand hiip(mh, mh, mh);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign qtqmqrax = qtqmqrax;
endmodule: zb

module mufdyip
  ( output wire logic [2:3][4:3]  lbvbtoneh
  , output wand logic [4:4] udhtsnmb [2:4][1:4][2:2][0:0]
  , output triand logic [4:2][3:0][1:4][1:3]  magkkejwv
  , input time fxoqmm [0:0][3:2][3:2]
  , input wire logic [2:2][2:1][2:3][1:2] n [2:4][3:2]
  , input tri0 logic [1:1][1:1][3:0][1:2] ncacylyp [4:1][2:4]
  , input tri logic [0:1] atjh [3:2][0:2]
  );
  
  
  xor hpdgl(lydrdoz, kp, lbvbtoneh);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> logic lbvbtoneh
  
  xor wdmhkmehe(kp, lbvbtoneh, lbvbtoneh);
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> logic lbvbtoneh
  //
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> logic lbvbtoneh
  
  nand xfvtt(bnxwqazlu, hc, dktaeu);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: mufdyip

module bvsg
  (output supply0 logic [3:3][2:2][3:3]  lt, output reg [2:3][2:1] httu [1:2]);
  
  wand logic [4:4] bjildsxhw [2:4][1:4][2:2][0:0];
  tri logic [0:1] yylkjprgt [3:2][0:2];
  tri0 logic [1:1][1:1][3:0][1:2] japryoybwc [4:1][2:4];
  wire logic [2:2][2:1][2:3][1:2] iubxhyizgz [2:4][3:2];
  time mc [0:0][3:2][3:2];
  
  not vnt(uk, ef);
  
  mufdyip gjb( .lbvbtoneh(gjz)
             , .udhtsnmb(bjildsxhw)
             , .magkkejwv(dsa)
             , .fxoqmm(mc)
             , .n(iubxhyizgz)
             , .ncacylyp(japryoybwc)
             , .atjh(yylkjprgt)
             );
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> wire logic gjz
  //
  // warning: implicit conversion of port connection truncates from 144 to 1 bits
  //   triand logic [4:2][3:0][1:4][1:3]  magkkejwv -> wire logic dsa
  
  not wkrq(gjz, krioulhy);
  
  
  // Single-driven assigns
  assign mc = '{'{'{'bz0,'bxz0},'{'bx1101,'b0x}}};
  assign httu = '{'{'{'b1,'b1x0},'{'b1zzz1,'bxxx}},'{'{'bz101,'b0z01},'{'bxz1x,'bzx}}};
  
  // Multi-driven assigns
  assign yylkjprgt = '{'{'{'b0xx,'b01001},'{'b0z,'b010z0},'{'b00,'b10}},'{'{'b010z,'bz0x},'{'bz1,'b1xz},'{'bx0,'b010x}}};
  assign iubxhyizgz = iubxhyizgz;
  assign uk = uk;
  assign japryoybwc = japryoybwc;
endmodule: bvsg

module zij
  ( output wand logic [4:4] ukpwknpeg [1:0][4:3][1:2][1:2]
  , output triand logic [2:3][0:0] hvebk [3:2][3:4][3:0]
  , output tri logic [4:2][0:3][4:3]  yzttip
  );
  
  wand logic [4:4] asd [2:4][1:4][2:2][0:0];
  wand logic [4:4] nkgor [2:4][1:4][2:2][0:0];
  reg [2:3][2:1] edxez [1:2];
  tri logic [0:1] ryns [3:2][0:2];
  tri0 logic [1:1][1:1][3:0][1:2] peod [4:1][2:4];
  time xtxlq [0:0][3:2][3:2];
  tri logic [0:1] ws [3:2][0:2];
  time myndlrfv [0:0][3:2][3:2];
  tri logic [0:1] cremgy [3:2][0:2];
  tri0 logic [1:1][1:1][3:0][1:2] zyos [4:1][2:4];
  wire logic [2:2][2:1][2:3][1:2] t [2:4][3:2];
  time xy [0:0][3:2][3:2];
  
  bvsg subxfa(.lt(ojjdfxwvwa), .httu(edxez));
  
  mufdyip tltemuos(.lbvbtoneh(gs), .udhtsnmb(nkgor), .magkkejwv(na), .fxoqmm(xy), .n(t), .ncacylyp(zyos), .atjh(cremgy));
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> wire logic gs
  //
  // warning: implicit conversion of port connection truncates from 144 to 1 bits
  //   triand logic [4:2][3:0][1:4][1:3]  magkkejwv -> wire logic na
  
  mufdyip jf(.lbvbtoneh(yzttip), .udhtsnmb(asd), .magkkejwv(qfuwag), .fxoqmm(myndlrfv), .n(t), .ncacylyp(zyos), .atjh(ws));
  // warning: implicit conversion of port connection expands from 4 to 24 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> tri logic [4:2][0:3][4:3]  yzttip
  //
  // warning: implicit conversion of port connection truncates from 144 to 1 bits
  //   triand logic [4:2][3:0][1:4][1:3]  magkkejwv -> wire logic qfuwag
  
  mufdyip eaxuk(.lbvbtoneh(gs), .udhtsnmb(nkgor), .magkkejwv(gs), .fxoqmm(xtxlq), .n(t), .ncacylyp(peod), .atjh(ryns));
  // warning: implicit conversion of port connection truncates from 4 to 1 bits
  //   wire logic [2:3][4:3]  lbvbtoneh -> wire logic gs
  //
  // warning: implicit conversion of port connection truncates from 144 to 1 bits
  //   triand logic [4:2][3:0][1:4][1:3]  magkkejwv -> wire logic gs
  
  
  // Single-driven assigns
  assign xtxlq = '{'{'{'b0z,'b0zx1},'{'bzz1,'bx}}};
  
  // Multi-driven assigns
  assign na = gs;
  assign peod = zyos;
  assign ryns = ws;
endmodule: zij



// Seed after: 10140135503795634854,5224943229413370507
