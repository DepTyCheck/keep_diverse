// Seed: 5024838802353150176,5224943229413370507

module vdazs
  ( output tri1 logic [1:2]  ywkj
  , output tri logic jirkjobk [3:3][0:0]
  , output bit xwq
  , output reg [0:4][1:4][2:4] bvy [3:2]
  , input supply0 logic [3:1][0:2][2:0][4:3] gxfxi [3:2][1:1][3:3]
  , input logic vhssam
  , input supply0 logic [4:2] iopfjros [0:0][4:1][0:4]
  , input logic tmo [3:2]
  );
  
  
  xor inrvwq(aa, ywkj, ywkj);
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri1 logic [1:2]  ywkj -> logic ywkj
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri1 logic [1:2]  ywkj -> logic ywkj
  
  not yrxnvcl(briy, vhssam);
  
  and jhykfst(xwq, ywkj, ywkj);
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic xwq -> bit xwq
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri1 logic [1:2]  ywkj -> logic ywkj
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  //   tri1 logic [1:2]  ywkj -> logic ywkj
  
  
  // Single-driven assigns
  assign bvy = bvy;
  
  // Multi-driven assigns
endmodule: vdazs

module vqfgruibl
  (output bit [2:0][3:4][4:2][0:3]  dbmkkcpyb, output bit h [2:0][3:3][2:2], output uwire logic [1:0][2:4] cyufnf [3:2][3:2]);
  
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: vqfgruibl

module eijyz
  (output trior logic [1:4][4:3][1:3] tlzajtwy [0:3][4:2][3:0], output logic [2:4][1:2] kmrxqr [2:0], output triand logic g);
  
  
  
  // Single-driven assigns
  assign kmrxqr = '{'{'{'b1z0,'b100},'{'bz10z,'b1xx},'{'bz0,'bx}},'{'{'b01z1,'b000},'{'b01x,'bzxx11},'{'b11z01,'b10zz}},'{'{'bx0,'b0x01},'{'b0x00x,'b1zzz},'{'b101z,'bx}}};
  
  // Multi-driven assigns
  assign tlzajtwy = tlzajtwy;
endmodule: eijyz



// Seed after: 14061539277969093024,5224943229413370507
