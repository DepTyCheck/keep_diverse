// Seed: 8288159748330704549,5224943229413370507

module fqzplwax
  ( output longint dvzhpk [2:3]
  , output uwire logic [4:2]  y
  , output supply1 logic [2:1][0:2]  zjgwfdylj
  , output wire logic [2:1][3:4][0:4][4:4] vr [4:3][0:3][4:3][0:1]
  );
  
  
  not zk(y, jqnhfadkbq);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  //   logic y -> uwire logic [4:2]  y
  
  not anuo(uo, xiseifukh);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign jqnhfadkbq = 'b1;
  assign xiseifukh = 'b10;
  assign vr = vr;
  assign zjgwfdylj = '{'{'bzz1z0,'b0110,'b1},'{'bx1x11,'bz11xz,'bz0x}};
endmodule: fqzplwax

module dpuimdbaza
  ( output tri0 logic gkkfdos [2:3][1:3]
  , output tri logic [1:1] tugqdj [0:3]
  , input triand logic vavhxnxf [1:2][0:0][3:3]
  , input bit [1:0] cdwdok [4:2][2:3]
  , input triand logic [4:4][4:1]  uekqsi
  , input uwire logic [2:0][2:2] ijckd [1:3]
  );
  
  
  or c(yco, vldb, vldb);
  
  not m(vldb, cjagsm);
  
  and djdvvugcv(bnv, vldb, bqvyzjq);
  
  not hnxvrjhq(jfengwj, fpe);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign tugqdj = tugqdj;
  assign gkkfdos = gkkfdos;
endmodule: dpuimdbaza

module pemitogpy
  ( output logic [4:4]  ysv
  , input tri0 logic [2:2][0:0][4:3][2:2] gmze [0:0]
  , input reg [3:4][4:2][0:4][2:4]  mpqncnvvl
  , input reg nr
  , input uwire logic khzpoghw [2:0][2:2]
  );
  
  
  and osma(chlznadxb, nr, nr);
  
  not a(chlznadxb, voxdp);
  
  not bagzzfqxj(enukqzcuj, voxdp);
  
  
  // Single-driven assigns
  assign ysv = ysv;
  
  // Multi-driven assigns
  assign voxdp = 'bz;
endmodule: pemitogpy



// Seed after: 4993766961193060316,5224943229413370507
