// Seed: 2232717311855488789,5224943229413370507

module vwaetrxxgw
  (output supply0 logic [1:0][2:1][1:0][2:1] ocw [0:0][1:1][0:0]);
  
  
  not psfwd(zcycypiey, e);
  
  xor euqd(mfabdcdwp, zcycypiey, nktfv);
  
  not jkmjs(e, jieclhy);
  
  not dpedk(nktfv, nktfv);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign mfabdcdwp = zcycypiey;
  assign jieclhy = 'b1111;
endmodule: vwaetrxxgw

module tmot
  ( output wor logic [3:3][3:2][2:3][4:3] yfwixz [0:4][1:0][3:4]
  , output bit [4:2]  fnzetuzm
  , output logic [2:1]  mnmwedlynr
  , input supply1 logic cif [0:3]
  , input reg dlwyfgp
  );
  
  supply0 logic [1:0][2:1][1:0][2:1] hv [0:0][1:1][0:0];
  
  vwaetrxxgw arbatytck(.ocw(hv));
  
  
  // Single-driven assigns
  assign fnzetuzm = fnzetuzm;
  assign mnmwedlynr = '{'b1z,'b1x};
  
  // Multi-driven assigns
endmodule: tmot



// Seed after: 12862203857658725940,5224943229413370507
