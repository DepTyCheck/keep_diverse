// Seed: 5678767469446421542,5224943229413370507

module a
  (output int namjubam, output uwire logic [2:1] eowh [3:3], input tri0 logic umuilwlv [4:4][3:0][3:3][2:3], input realtime o);
  
  
  nand lksvhqytmg(namjubam, namjubam, namjubam);
  // warning: implicit conversion of port connection expands from 1 to 32 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic namjubam -> int namjubam
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int namjubam -> logic namjubam
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int namjubam -> logic namjubam
  
  not drzmvldm(dscwczc, o);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime o -> logic o
  
  
  // Single-driven assigns
  assign eowh = eowh;
  
  // Multi-driven assigns
endmodule: a

module jsnjwosnhh
  ( output triand logic [2:2][1:0][2:4] tpwlrk [1:1][3:2][1:2][1:3]
  , output shortint fvjwvuvf
  , output logic [0:4][3:4]  uueap
  , output wor logic [0:2] fiknw [3:0]
  , input logic rnd
  , input wand logic [2:1] dz [1:1][3:1][1:2][0:2]
  , input triand logic [1:3][0:4] ozo [2:4][1:0][0:4]
  , input reg [4:3][1:1]  ccxs
  );
  
  
  
  // Single-driven assigns
  assign uueap = '{'{'bxz1,'bzx},'{'bx0z,'b001},'{'bzz1,'bx0xx0},'{'bx0011,'b0zx0},'{'b0x,'b000xz}};
  assign fvjwvuvf = fvjwvuvf;
  
  // Multi-driven assigns
  assign tpwlrk = tpwlrk;
  assign fiknw = '{'{'b0zz1,'b0xz,'bxz},'{'b0zx,'bx,'b0x},'{'bx01xz,'b11,'bx},'{'b1zzx0,'bz1x10,'bz}};
endmodule: jsnjwosnhh

module fwll
  ( output time fzbybdnbmt
  , output real uhrymn
  , output wor logic slmvvprj [0:1][2:4]
  , input reg [0:3][0:2][3:3] go [2:0]
  , input shortreal sh
  );
  
  uwire logic [2:1] xyfqtrzng [3:3];
  tri0 logic sokftyjtd [4:4][3:0][3:3][2:3];
  
  a jboyrclh(.namjubam(fqkqasi), .eowh(xyfqtrzng), .umuilwlv(sokftyjtd), .o(fzbybdnbmt));
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int namjubam -> wire logic fqkqasi
  //
  // warning: implicit conversion changes signedness from unsigned to signed
  //   time fzbybdnbmt -> realtime o
  
  and jkoqig(fzbybdnbmt, ykhlhxlhsh, md);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  //   logic fzbybdnbmt -> time fzbybdnbmt
  
  or zbqzwmpn(el, fzbybdnbmt, ykhlhxlhsh);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  //   time fzbybdnbmt -> logic fzbybdnbmt
  
  
  // Single-driven assigns
  assign uhrymn = fqkqasi;
  
  // Multi-driven assigns
endmodule: fwll



// Seed after: 10034344404040501477,5224943229413370507
