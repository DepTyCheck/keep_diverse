// Seed: 16723051014337592514,5224943229413370507

module swhgfquum
  (output supply0 logic yrjc [3:3], input tri logic [3:2] okxembmzrz [2:1][2:0][2:0][0:4], input supply1 logic iclxy [1:0]);
  
  
  xor yuzprfweh(whtajdd, jj, jj);
  
  nand bsf(e, whtajdd, efdx);
  
  nand qyn(e, jj, aqcsxi);
  
  nand enpcaive(e, jqchiosoka, obz);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign jqchiosoka = whtajdd;
  assign yrjc = '{'bz1};
  assign jj = 'bzzz;
endmodule: swhgfquum



// Seed after: 12436611882516698977,5224943229413370507
