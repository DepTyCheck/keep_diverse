// Seed: 7718581316640303111,5224943229413370507

module pxvth
  ( output supply1 logic x
  , output logic [2:0][2:1][4:4][1:0]  hufuakrxu
  , output bit [4:3][4:4][3:0][1:1]  mvqymitgli
  , input supply1 logic [2:1][2:3][0:2][0:4]  gropup
  , input uwire logic [0:3] wal [2:3][2:2]
  , input tri0 logic [3:1][3:2][1:4] gpco [3:4]
  );
  
  
  not azoxr(ne, jvq);
  
  xor axankmfqa(wqkweu, mvqymitgli, lchrousw);
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:3][4:4][3:0][1:1]  mvqymitgli -> logic mvqymitgli
  
  xor atv(hufuakrxu, x, ejinoanh);
  // warning: implicit conversion of port connection expands from 1 to 12 bits
  //   logic hufuakrxu -> logic [2:0][2:1][4:4][1:0]  hufuakrxu
  
  
  // Single-driven assigns
  assign mvqymitgli = x;
  
  // Multi-driven assigns
endmodule: pxvth

module dlefkpbl
  (output tri0 logic htig [2:3][0:0][0:1][2:2], output realtime nwqtvajbci);
  
  tri0 logic [3:1][3:2][1:4] stgl [3:4];
  uwire logic [0:3] vnhefpilbx [2:3][2:2];
  
  not wsucooma(nwqtvajbci, nwqtvajbci);
  // warning: implicit conversion of port connection expands from 1 to 64 bits
  // warning: implicit conversion changes signedness from unsigned to signed
  //   logic nwqtvajbci -> realtime nwqtvajbci
  //
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime nwqtvajbci -> logic nwqtvajbci
  
  nand ydavjtk(ch, cwdt, nwqtvajbci);
  // warning: implicit conversion of port connection truncates from 64 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime nwqtvajbci -> logic nwqtvajbci
  
  not tbbu(cwdt, tne);
  
  pxvth ledlmd(.x(uqtnws), .hufuakrxu(yncihbw), .mvqymitgli(byiyzqayln), .gropup(nwqtvajbci), .wal(vnhefpilbx), .gpco(stgl));
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [2:0][2:1][4:4][1:0]  hufuakrxu -> wire logic yncihbw
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [4:3][4:4][3:0][1:1]  mvqymitgli -> wire logic byiyzqayln
  //
  // warning: implicit conversion of port connection truncates from 64 to 60 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   realtime nwqtvajbci -> supply1 logic [2:1][2:3][0:2][0:4]  gropup
  
  
  // Single-driven assigns
  assign vnhefpilbx = '{'{'{'b0xzz,'b1x0,'bz0,'bzzxzz}},'{'{'bz,'b000,'b11z1,'b1z}}};
  
  // Multi-driven assigns
endmodule: dlefkpbl

module ojrn
  (output tri1 logic [2:1][1:3][2:0]  ww, input supply0 logic wez [0:4][3:1][2:3], input wand logic [1:4][0:3][4:4] jhv [0:0]);
  
  
  xor cgixteammt(oc, coxx, ltsjvkn);
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign ltsjvkn = ww;
  assign coxx = ww;
endmodule: ojrn



// Seed after: 7587504049292560125,5224943229413370507
