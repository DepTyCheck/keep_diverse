// Seed: 4214566392895304490,5224943229413370507

module xtwipi
  (output wire logic duo [3:2][0:3], output wor logic tsuy [3:4], input bit [0:0][2:0][0:2]  ucbjrmed);
  
  
  and gcgaaoc(ibcjnah, ucbjrmed, ucbjrmed);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:0][2:0][0:2]  ucbjrmed -> logic ucbjrmed
  //
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:0][2:0][0:2]  ucbjrmed -> logic ucbjrmed
  
  nand vamejkrj(ibcjnah, ucbjrmed, ibcjnah);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:0][2:0][0:2]  ucbjrmed -> logic ucbjrmed
  
  nand uvinq(cgvfifsyw, cgvfifsyw, ibcjnah);
  
  not nbelqumvd(ibcjnah, ucbjrmed);
  // warning: implicit conversion of port connection truncates from 9 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [0:0][2:0][0:2]  ucbjrmed -> logic ucbjrmed
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign duo = '{'{'bx11x,'bz,'b0z,'b0z0zx},'{'bx,'b0xz0,'b00,'bz1zz}};
  assign tsuy = tsuy;
endmodule: xtwipi

module y
  ( output tri1 logic [0:1][0:0][1:3] dxwsl [4:2]
  , output logic wlcgz [1:3][3:4]
  , output tri1 logic [0:1][3:2][3:2][2:3]  oh
  , input triand logic [0:0] sqnpddyno [3:1][2:0][4:2][2:4]
  , input shortreal eqqrcihajj
  );
  
  
  xor mtmgctgi(tpjgpokryi, eqqrcihajj, oh);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal eqqrcihajj -> logic eqqrcihajj
  //
  // warning: implicit conversion of port connection truncates from 16 to 1 bits
  //   tri1 logic [0:1][3:2][3:2][2:3]  oh -> logic oh
  
  nand ke(oh, lvmvx, abfgmr);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  //   logic oh -> tri1 logic [0:1][3:2][3:2][2:3]  oh
  
  not sf(oh, koujrqmgvi);
  // warning: implicit conversion of port connection expands from 1 to 16 bits
  //   logic oh -> tri1 logic [0:1][3:2][3:2][2:3]  oh
  
  nand ftdogecops(ksl, eqqrcihajj, cxdnqlmz);
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  //   shortreal eqqrcihajj -> logic eqqrcihajj
  
  
  // Single-driven assigns
  assign wlcgz = '{'{'b01zxx,'b0x},'{'b0xx1,'bx},'{'bx0xx,'bxx}};
  
  // Multi-driven assigns
  assign koujrqmgvi = 'b0zz;
endmodule: y



// Seed after: 31107661655320341,5224943229413370507
