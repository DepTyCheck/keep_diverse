// Seed: 13115324323945111150,5224943229413370507

module tztnwfbby
  (input tri logic [3:3][2:0][1:2][0:3]  kl, input logic [1:0][3:1][3:2]  otcfcybf, input reg [2:3][1:2][3:0][2:3]  souaft);
  
  
  not dl(kl, kl);
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   logic kl -> tri logic [3:3][2:0][1:2][0:3]  kl
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   tri logic [3:3][2:0][1:2][0:3]  kl -> logic kl
  
  xor plb(kl, kl, kl);
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   logic kl -> tri logic [3:3][2:0][1:2][0:3]  kl
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   tri logic [3:3][2:0][1:2][0:3]  kl -> logic kl
  //
  // warning: implicit conversion of port connection truncates from 24 to 1 bits
  //   tri logic [3:3][2:0][1:2][0:3]  kl -> logic kl
  
  and aaihohgo(kl, otcfcybf, souaft);
  // warning: implicit conversion of port connection expands from 1 to 24 bits
  //   logic kl -> tri logic [3:3][2:0][1:2][0:3]  kl
  //
  // warning: implicit conversion of port connection truncates from 12 to 1 bits
  //   logic [1:0][3:1][3:2]  otcfcybf -> logic otcfcybf
  //
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  //   reg [2:3][1:2][3:0][2:3]  souaft -> logic souaft
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
  assign kl = '{'{'{'{'bx1,'b00,'bx00,'bx},'{'b00x1,'bzz0z,'b0zx,'bz10z}},'{'{'b0x0,'b1xx,'bzz,'bx0z0x},'{'b0zz0z,'bx,'b00,'b0z1x}},'{'{'b1z0x,'b1,'b0,'b10},'{'b0z01,'b01,'b1xz,'b111z}}}};
endmodule: tztnwfbby

module ltadt
  (output bit [2:4]  mufdoz, input reg [0:4][1:2][4:3] ky [4:4], input reg [2:4][1:2][4:1] rhylpfrnri [2:2], input byte uiktpzfmgu);
  
  
  not hguwtzxzfd(rpibz, mufdoz);
  // warning: implicit conversion of port connection truncates from 3 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:4]  mufdoz -> logic mufdoz
  
  and ng(mufdoz, uiktpzfmgu, szirszuzt);
  // warning: implicit conversion of port connection expands from 1 to 3 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic mufdoz -> bit [2:4]  mufdoz
  //
  // warning: implicit conversion of port connection truncates from 8 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   byte uiktpzfmgu -> logic uiktpzfmgu
  
  
  // Single-driven assigns
  
  // Multi-driven assigns
endmodule: ltadt



// Seed after: 12435502455885098234,5224943229413370507
